module compressor(
      input wire [63:0] src00,
      input wire [63:0] src01,
      input wire [63:0] src02,
      input wire [63:0] src03,
      input wire [63:0] src04,
      input wire [63:0] src05,
      input wire [63:0] src06,
      input wire [63:0] src07,
      input wire [63:0] src08,
      input wire [63:0] src09,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      input wire [63:0] src32,
      input wire [63:0] src33,
      input wire [63:0] src34,
      input wire [63:0] src35,
      input wire [63:0] src36,
      input wire [63:0] src37,
      input wire [63:0] src38,
      input wire [63:0] src39,
      input wire [63:0] src40,
      input wire [63:0] src41,
      input wire [63:0] src42,
      input wire [63:0] src43,
      input wire [63:0] src44,
      input wire [63:0] src45,
      input wire [63:0] src46,
      input wire [63:0] src47,
      input wire [63:0] src48,
      input wire [63:0] src49,
      input wire [63:0] src50,
      input wire [63:0] src51,
      input wire [63:0] src52,
      input wire [63:0] src53,
      input wire [63:0] src54,
      input wire [63:0] src55,
      input wire [63:0] src56,
      input wire [63:0] src57,
      input wire [63:0] src58,
      input wire [63:0] src59,
      input wire [63:0] src60,
      input wire [63:0] src61,
      input wire [63:0] src62,
      input wire [63:0] src63,
      output wire [1:0] dst00,
      output wire [0:0] dst01,
      output wire [1:0] dst02,
      output wire [1:0] dst03,
      output wire [1:0] dst04,
      output wire [1:0] dst05,
      output wire [1:0] dst06,
      output wire [1:0] dst07,
      output wire [0:0] dst08,
      output wire [1:0] dst09,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [0:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [0:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [0:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [0:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [0:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [0:0] dst70
   );
   wire [101:0] stage00;
   wire [130:0] stage01;
   wire [120:0] stage02;
   wire [142:0] stage03;
   wire [127:0] stage04;
   wire [131:0] stage05;
   wire [122:0] stage06;
   wire [123:0] stage07;
   wire [129:0] stage08;
   wire [177:0] stage09;
   wire [148:0] stage10;
   wire [161:0] stage11;
   wire [157:0] stage12;
   wire [143:0] stage13;
   wire [120:0] stage14;
   wire [172:0] stage15;
   wire [117:0] stage16;
   wire [160:0] stage17;
   wire [131:0] stage18;
   wire [136:0] stage19;
   wire [157:0] stage20;
   wire [121:0] stage21;
   wire [126:0] stage22;
   wire [149:0] stage23;
   wire [127:0] stage24;
   wire [140:0] stage25;
   wire [118:0] stage26;
   wire [151:0] stage27;
   wire [151:0] stage28;
   wire [118:0] stage29;
   wire [138:0] stage30;
   wire [129:0] stage31;
   wire [117:0] stage32;
   wire [116:0] stage33;
   wire [123:0] stage34;
   wire [117:0] stage35;
   wire [150:0] stage36;
   wire [130:0] stage37;
   wire [122:0] stage38;
   wire [120:0] stage39;
   wire [144:0] stage40;
   wire [148:0] stage41;
   wire [144:0] stage42;
   wire [160:0] stage43;
   wire [129:0] stage44;
   wire [143:0] stage45;
   wire [136:0] stage46;
   wire [138:0] stage47;
   wire [131:0] stage48;
   wire [153:0] stage49;
   wire [126:0] stage50;
   wire [121:0] stage51;
   wire [123:0] stage52;
   wire [126:0] stage53;
   wire [140:0] stage54;
   wire [118:0] stage55;
   wire [156:0] stage56;
   wire [129:0] stage57;
   wire [127:0] stage58;
   wire [145:0] stage59;
   wire [139:0] stage60;
   wire [151:0] stage61;
   wire [137:0] stage62;
   wire [121:0] stage63;
   wire [51:0] stage64;
   wire [38:0] stage65;
   wire [16:0] stage66;
   wire [8:0] stage67;
   wire [3:0] stage68;
   wire [2:0] stage69;
   wire [0:0] stage70;
   assign stage00[63:0] = src00;
   assign stage01[63:0] = src01;
   assign stage02[63:0] = src02;
   assign stage03[63:0] = src03;
   assign stage04[63:0] = src04;
   assign stage05[63:0] = src05;
   assign stage06[63:0] = src06;
   assign stage07[63:0] = src07;
   assign stage08[63:0] = src08;
   assign stage09[63:0] = src09;
   assign stage10[63:0] = src10;
   assign stage11[63:0] = src11;
   assign stage12[63:0] = src12;
   assign stage13[63:0] = src13;
   assign stage14[63:0] = src14;
   assign stage15[63:0] = src15;
   assign stage16[63:0] = src16;
   assign stage17[63:0] = src17;
   assign stage18[63:0] = src18;
   assign stage19[63:0] = src19;
   assign stage20[63:0] = src20;
   assign stage21[63:0] = src21;
   assign stage22[63:0] = src22;
   assign stage23[63:0] = src23;
   assign stage24[63:0] = src24;
   assign stage25[63:0] = src25;
   assign stage26[63:0] = src26;
   assign stage27[63:0] = src27;
   assign stage28[63:0] = src28;
   assign stage29[63:0] = src29;
   assign stage30[63:0] = src30;
   assign stage31[63:0] = src31;
   assign stage32[63:0] = src32;
   assign stage33[63:0] = src33;
   assign stage34[63:0] = src34;
   assign stage35[63:0] = src35;
   assign stage36[63:0] = src36;
   assign stage37[63:0] = src37;
   assign stage38[63:0] = src38;
   assign stage39[63:0] = src39;
   assign stage40[63:0] = src40;
   assign stage41[63:0] = src41;
   assign stage42[63:0] = src42;
   assign stage43[63:0] = src43;
   assign stage44[63:0] = src44;
   assign stage45[63:0] = src45;
   assign stage46[63:0] = src46;
   assign stage47[63:0] = src47;
   assign stage48[63:0] = src48;
   assign stage49[63:0] = src49;
   assign stage50[63:0] = src50;
   assign stage51[63:0] = src51;
   assign stage52[63:0] = src52;
   assign stage53[63:0] = src53;
   assign stage54[63:0] = src54;
   assign stage55[63:0] = src55;
   assign stage56[63:0] = src56;
   assign stage57[63:0] = src57;
   assign stage58[63:0] = src58;
   assign stage59[63:0] = src59;
   assign stage60[63:0] = src60;
   assign stage61[63:0] = src61;
   assign stage62[63:0] = src62;
   assign stage63[63:0] = src63;
   assign dst00 = stage00[101:100];
   assign dst01 = stage01[130:130];
   assign dst02 = stage02[120:119];
   assign dst03 = stage03[142:141];
   assign dst04 = stage04[127:126];
   assign dst05 = stage05[131:130];
   assign dst06 = stage06[122:121];
   assign dst07 = stage07[123:122];
   assign dst08 = stage08[129:129];
   assign dst09 = stage09[177:176];
   assign dst10 = stage10[148:147];
   assign dst11 = stage11[161:160];
   assign dst12 = stage12[157:156];
   assign dst13 = stage13[143:142];
   assign dst14 = stage14[120:119];
   assign dst15 = stage15[172:171];
   assign dst16 = stage16[117:116];
   assign dst17 = stage17[160:159];
   assign dst18 = stage18[131:130];
   assign dst19 = stage19[136:135];
   assign dst20 = stage20[157:157];
   assign dst21 = stage21[121:120];
   assign dst22 = stage22[126:125];
   assign dst23 = stage23[149:148];
   assign dst24 = stage24[127:126];
   assign dst25 = stage25[140:139];
   assign dst26 = stage26[118:117];
   assign dst27 = stage27[151:150];
   assign dst28 = stage28[151:150];
   assign dst29 = stage29[118:117];
   assign dst30 = stage30[138:137];
   assign dst31 = stage31[129:129];
   assign dst32 = stage32[117:116];
   assign dst33 = stage33[116:115];
   assign dst34 = stage34[123:123];
   assign dst35 = stage35[117:116];
   assign dst36 = stage36[150:149];
   assign dst37 = stage37[130:129];
   assign dst38 = stage38[122:121];
   assign dst39 = stage39[120:119];
   assign dst40 = stage40[144:143];
   assign dst41 = stage41[148:147];
   assign dst42 = stage42[144:143];
   assign dst43 = stage43[160:159];
   assign dst44 = stage44[129:128];
   assign dst45 = stage45[143:142];
   assign dst46 = stage46[136:136];
   assign dst47 = stage47[138:137];
   assign dst48 = stage48[131:130];
   assign dst49 = stage49[153:152];
   assign dst50 = stage50[126:125];
   assign dst51 = stage51[121:120];
   assign dst52 = stage52[123:122];
   assign dst53 = stage53[126:125];
   assign dst54 = stage54[140:139];
   assign dst55 = stage55[118:117];
   assign dst56 = stage56[156:155];
   assign dst57 = stage57[129:128];
   assign dst58 = stage58[127:127];
   assign dst59 = stage59[145:144];
   assign dst60 = stage60[139:138];
   assign dst61 = stage61[151:150];
   assign dst62 = stage62[137:136];
   assign dst63 = stage63[121:120];
   assign dst64 = stage64[51:51];
   assign dst65 = stage65[38:37];
   assign dst66 = stage66[16:15];
   assign dst67 = stage67[8:7];
   assign dst68 = stage68[3:2];
   assign dst69 = stage69[2:1];
   assign dst70 = stage70[0:0];
   gpc1_1 gpc1_1_0(
      {stage00[0]},
      {stage00[64]}
   );
   gpc1_1 gpc1_1_1(
      {stage00[1]},
      {stage00[65]}
   );
   gpc1_1 gpc1_1_2(
      {stage00[2]},
      {stage00[66]}
   );
   gpc1_1 gpc1_1_3(
      {stage00[3]},
      {stage00[67]}
   );
   gpc615_5 gpc615_5_4(
      {stage00[4], stage00[5], stage00[6], stage00[7], stage00[8]},
      {stage01[0]},
      {stage02[0], stage02[1], stage02[2], stage02[3], stage02[4], stage02[5]},
      {stage04[64], stage03[64], stage02[64], stage01[64], stage00[68]}
   );
   gpc615_5 gpc615_5_5(
      {stage00[9], stage00[10], stage00[11], stage00[12], stage00[13]},
      {stage01[1]},
      {stage02[6], stage02[7], stage02[8], stage02[9], stage02[10], stage02[11]},
      {stage04[65], stage03[65], stage02[65], stage01[65], stage00[69]}
   );
   gpc615_5 gpc615_5_6(
      {stage00[14], stage00[15], stage00[16], stage00[17], stage00[18]},
      {stage01[2]},
      {stage02[12], stage02[13], stage02[14], stage02[15], stage02[16], stage02[17]},
      {stage04[66], stage03[66], stage02[66], stage01[66], stage00[70]}
   );
   gpc615_5 gpc615_5_7(
      {stage00[19], stage00[20], stage00[21], stage00[22], stage00[23]},
      {stage01[3]},
      {stage02[18], stage02[19], stage02[20], stage02[21], stage02[22], stage02[23]},
      {stage04[67], stage03[67], stage02[67], stage01[67], stage00[71]}
   );
   gpc615_5 gpc615_5_8(
      {stage00[24], stage00[25], stage00[26], stage00[27], stage00[28]},
      {stage01[4]},
      {stage02[24], stage02[25], stage02[26], stage02[27], stage02[28], stage02[29]},
      {stage04[68], stage03[68], stage02[68], stage01[68], stage00[72]}
   );
   gpc2135_5 gpc2135_5_9(
      {stage00[29], stage00[30], stage00[31], stage00[32], stage00[33]},
      {stage01[5], stage01[6], stage01[7]},
      {stage02[30]},
      {stage03[0], stage03[1]},
      {stage04[69], stage03[69], stage02[69], stage01[69], stage00[73]}
   );
   gpc2135_5 gpc2135_5_10(
      {stage00[34], stage00[35], stage00[36], stage00[37], stage00[38]},
      {stage01[8], stage01[9], stage01[10]},
      {stage02[31]},
      {stage03[2], stage03[3]},
      {stage04[70], stage03[70], stage02[70], stage01[70], stage00[74]}
   );
   gpc2135_5 gpc2135_5_11(
      {stage00[39], stage00[40], stage00[41], stage00[42], stage00[43]},
      {stage01[11], stage01[12], stage01[13]},
      {stage02[32]},
      {stage03[4], stage03[5]},
      {stage04[71], stage03[71], stage02[71], stage01[71], stage00[75]}
   );
   gpc2135_5 gpc2135_5_12(
      {stage00[44], stage00[45], stage00[46], stage00[47], stage00[48]},
      {stage01[14], stage01[15], stage01[16]},
      {stage02[33]},
      {stage03[6], stage03[7]},
      {stage04[72], stage03[72], stage02[72], stage01[72], stage00[76]}
   );
   gpc2135_5 gpc2135_5_13(
      {stage00[49], stage00[50], stage00[51], stage00[52], stage00[53]},
      {stage01[17], stage01[18], stage01[19]},
      {stage02[34]},
      {stage03[8], stage03[9]},
      {stage04[73], stage03[73], stage02[73], stage01[73], stage00[77]}
   );
   gpc2135_5 gpc2135_5_14(
      {stage00[54], stage00[55], stage00[56], stage00[57], stage00[58]},
      {stage01[20], stage01[21], stage01[22]},
      {stage02[35]},
      {stage03[10], stage03[11]},
      {stage04[74], stage03[74], stage02[74], stage01[74], stage00[78]}
   );
   gpc2135_5 gpc2135_5_15(
      {stage00[59], stage00[60], stage00[61], stage00[62], stage00[63]},
      {stage01[23], stage01[24], stage01[25]},
      {stage02[36]},
      {stage03[12], stage03[13]},
      {stage04[75], stage03[75], stage02[75], stage01[75], stage00[79]}
   );
   gpc1_1 gpc1_1_16(
      {stage01[26]},
      {stage01[76]}
   );
   gpc1_1 gpc1_1_17(
      {stage01[27]},
      {stage01[77]}
   );
   gpc1_1 gpc1_1_18(
      {stage01[28]},
      {stage01[78]}
   );
   gpc1_1 gpc1_1_19(
      {stage01[29]},
      {stage01[79]}
   );
   gpc1_1 gpc1_1_20(
      {stage01[30]},
      {stage01[80]}
   );
   gpc1_1 gpc1_1_21(
      {stage01[31]},
      {stage01[81]}
   );
   gpc1_1 gpc1_1_22(
      {stage01[32]},
      {stage01[82]}
   );
   gpc1_1 gpc1_1_23(
      {stage01[33]},
      {stage01[83]}
   );
   gpc1_1 gpc1_1_24(
      {stage01[34]},
      {stage01[84]}
   );
   gpc1_1 gpc1_1_25(
      {stage01[35]},
      {stage01[85]}
   );
   gpc1_1 gpc1_1_26(
      {stage01[36]},
      {stage01[86]}
   );
   gpc1_1 gpc1_1_27(
      {stage01[37]},
      {stage01[87]}
   );
   gpc1_1 gpc1_1_28(
      {stage01[38]},
      {stage01[88]}
   );
   gpc1_1 gpc1_1_29(
      {stage01[39]},
      {stage01[89]}
   );
   gpc1_1 gpc1_1_30(
      {stage01[40]},
      {stage01[90]}
   );
   gpc1_1 gpc1_1_31(
      {stage01[41]},
      {stage01[91]}
   );
   gpc1_1 gpc1_1_32(
      {stage01[42]},
      {stage01[92]}
   );
   gpc1_1 gpc1_1_33(
      {stage01[43]},
      {stage01[93]}
   );
   gpc1_1 gpc1_1_34(
      {stage01[44]},
      {stage01[94]}
   );
   gpc1_1 gpc1_1_35(
      {stage01[45]},
      {stage01[95]}
   );
   gpc1_1 gpc1_1_36(
      {stage01[46]},
      {stage01[96]}
   );
   gpc1_1 gpc1_1_37(
      {stage01[47]},
      {stage01[97]}
   );
   gpc1_1 gpc1_1_38(
      {stage01[48]},
      {stage01[98]}
   );
   gpc1_1 gpc1_1_39(
      {stage01[49]},
      {stage01[99]}
   );
   gpc1_1 gpc1_1_40(
      {stage01[50]},
      {stage01[100]}
   );
   gpc1_1 gpc1_1_41(
      {stage01[51]},
      {stage01[101]}
   );
   gpc1_1 gpc1_1_42(
      {stage01[52]},
      {stage01[102]}
   );
   gpc1_1 gpc1_1_43(
      {stage01[53]},
      {stage01[103]}
   );
   gpc1_1 gpc1_1_44(
      {stage01[54]},
      {stage01[104]}
   );
   gpc1_1 gpc1_1_45(
      {stage01[55]},
      {stage01[105]}
   );
   gpc1_1 gpc1_1_46(
      {stage01[56]},
      {stage01[106]}
   );
   gpc1_1 gpc1_1_47(
      {stage01[57]},
      {stage01[107]}
   );
   gpc1_1 gpc1_1_48(
      {stage01[58]},
      {stage01[108]}
   );
   gpc2135_5 gpc2135_5_49(
      {stage01[59], stage01[60], stage01[61], stage01[62], stage01[63]},
      {stage02[37], stage02[38], stage02[39]},
      {stage03[14]},
      {stage04[0], stage04[1]},
      {stage05[64], stage04[76], stage03[76], stage02[76], stage01[109]}
   );
   gpc1_1 gpc1_1_50(
      {stage02[40]},
      {stage02[77]}
   );
   gpc1_1 gpc1_1_51(
      {stage02[41]},
      {stage02[78]}
   );
   gpc1_1 gpc1_1_52(
      {stage02[42]},
      {stage02[79]}
   );
   gpc1_1 gpc1_1_53(
      {stage02[43]},
      {stage02[80]}
   );
   gpc1_1 gpc1_1_54(
      {stage02[44]},
      {stage02[81]}
   );
   gpc1_1 gpc1_1_55(
      {stage02[45]},
      {stage02[82]}
   );
   gpc606_5 gpc606_5_56(
      {stage02[46], stage02[47], stage02[48], stage02[49], stage02[50], stage02[51]},
      {stage04[2], stage04[3], stage04[4], stage04[5], stage04[6], stage04[7]},
      {stage06[64], stage05[65], stage04[77], stage03[77], stage02[83]}
   );
   gpc606_5 gpc606_5_57(
      {stage02[52], stage02[53], stage02[54], stage02[55], stage02[56], stage02[57]},
      {stage04[8], stage04[9], stage04[10], stage04[11], stage04[12], stage04[13]},
      {stage06[65], stage05[66], stage04[78], stage03[78], stage02[84]}
   );
   gpc606_5 gpc606_5_58(
      {stage02[58], stage02[59], stage02[60], stage02[61], stage02[62], stage02[63]},
      {stage04[14], stage04[15], stage04[16], stage04[17], stage04[18], stage04[19]},
      {stage06[66], stage05[67], stage04[79], stage03[79], stage02[85]}
   );
   gpc1_1 gpc1_1_59(
      {stage03[15]},
      {stage03[80]}
   );
   gpc1_1 gpc1_1_60(
      {stage03[16]},
      {stage03[81]}
   );
   gpc1_1 gpc1_1_61(
      {stage03[17]},
      {stage03[82]}
   );
   gpc1_1 gpc1_1_62(
      {stage03[18]},
      {stage03[83]}
   );
   gpc1_1 gpc1_1_63(
      {stage03[19]},
      {stage03[84]}
   );
   gpc1_1 gpc1_1_64(
      {stage03[20]},
      {stage03[85]}
   );
   gpc1_1 gpc1_1_65(
      {stage03[21]},
      {stage03[86]}
   );
   gpc1_1 gpc1_1_66(
      {stage03[22]},
      {stage03[87]}
   );
   gpc1_1 gpc1_1_67(
      {stage03[23]},
      {stage03[88]}
   );
   gpc1_1 gpc1_1_68(
      {stage03[24]},
      {stage03[89]}
   );
   gpc1_1 gpc1_1_69(
      {stage03[25]},
      {stage03[90]}
   );
   gpc1_1 gpc1_1_70(
      {stage03[26]},
      {stage03[91]}
   );
   gpc1_1 gpc1_1_71(
      {stage03[27]},
      {stage03[92]}
   );
   gpc1_1 gpc1_1_72(
      {stage03[28]},
      {stage03[93]}
   );
   gpc1_1 gpc1_1_73(
      {stage03[29]},
      {stage03[94]}
   );
   gpc1_1 gpc1_1_74(
      {stage03[30]},
      {stage03[95]}
   );
   gpc1_1 gpc1_1_75(
      {stage03[31]},
      {stage03[96]}
   );
   gpc1_1 gpc1_1_76(
      {stage03[32]},
      {stage03[97]}
   );
   gpc1_1 gpc1_1_77(
      {stage03[33]},
      {stage03[98]}
   );
   gpc1_1 gpc1_1_78(
      {stage03[34]},
      {stage03[99]}
   );
   gpc1_1 gpc1_1_79(
      {stage03[35]},
      {stage03[100]}
   );
   gpc1_1 gpc1_1_80(
      {stage03[36]},
      {stage03[101]}
   );
   gpc1_1 gpc1_1_81(
      {stage03[37]},
      {stage03[102]}
   );
   gpc1_1 gpc1_1_82(
      {stage03[38]},
      {stage03[103]}
   );
   gpc1_1 gpc1_1_83(
      {stage03[39]},
      {stage03[104]}
   );
   gpc1_1 gpc1_1_84(
      {stage03[40]},
      {stage03[105]}
   );
   gpc1_1 gpc1_1_85(
      {stage03[41]},
      {stage03[106]}
   );
   gpc1_1 gpc1_1_86(
      {stage03[42]},
      {stage03[107]}
   );
   gpc1_1 gpc1_1_87(
      {stage03[43]},
      {stage03[108]}
   );
   gpc1_1 gpc1_1_88(
      {stage03[44]},
      {stage03[109]}
   );
   gpc1_1 gpc1_1_89(
      {stage03[45]},
      {stage03[110]}
   );
   gpc1_1 gpc1_1_90(
      {stage03[46]},
      {stage03[111]}
   );
   gpc1_1 gpc1_1_91(
      {stage03[47]},
      {stage03[112]}
   );
   gpc1_1 gpc1_1_92(
      {stage03[48]},
      {stage03[113]}
   );
   gpc1_1 gpc1_1_93(
      {stage03[49]},
      {stage03[114]}
   );
   gpc1_1 gpc1_1_94(
      {stage03[50]},
      {stage03[115]}
   );
   gpc1_1 gpc1_1_95(
      {stage03[51]},
      {stage03[116]}
   );
   gpc1_1 gpc1_1_96(
      {stage03[52]},
      {stage03[117]}
   );
   gpc1_1 gpc1_1_97(
      {stage03[53]},
      {stage03[118]}
   );
   gpc615_5 gpc615_5_98(
      {stage03[54], stage03[55], stage03[56], stage03[57], stage03[58]},
      {stage04[20]},
      {stage05[0], stage05[1], stage05[2], stage05[3], stage05[4], stage05[5]},
      {stage07[64], stage06[67], stage05[68], stage04[80], stage03[119]}
   );
   gpc615_5 gpc615_5_99(
      {stage03[59], stage03[60], stage03[61], stage03[62], stage03[63]},
      {stage04[21]},
      {stage05[6], stage05[7], stage05[8], stage05[9], stage05[10], stage05[11]},
      {stage07[65], stage06[68], stage05[69], stage04[81], stage03[120]}
   );
   gpc1_1 gpc1_1_100(
      {stage04[22]},
      {stage04[82]}
   );
   gpc1_1 gpc1_1_101(
      {stage04[23]},
      {stage04[83]}
   );
   gpc1_1 gpc1_1_102(
      {stage04[24]},
      {stage04[84]}
   );
   gpc1_1 gpc1_1_103(
      {stage04[25]},
      {stage04[85]}
   );
   gpc606_5 gpc606_5_104(
      {stage04[26], stage04[27], stage04[28], stage04[29], stage04[30], stage04[31]},
      {stage06[0], stage06[1], stage06[2], stage06[3], stage06[4], stage06[5]},
      {stage08[64], stage07[66], stage06[69], stage05[70], stage04[86]}
   );
   gpc606_5 gpc606_5_105(
      {stage04[32], stage04[33], stage04[34], stage04[35], stage04[36], stage04[37]},
      {stage06[6], stage06[7], stage06[8], stage06[9], stage06[10], stage06[11]},
      {stage08[65], stage07[67], stage06[70], stage05[71], stage04[87]}
   );
   gpc606_5 gpc606_5_106(
      {stage04[38], stage04[39], stage04[40], stage04[41], stage04[42], stage04[43]},
      {stage06[12], stage06[13], stage06[14], stage06[15], stage06[16], stage06[17]},
      {stage08[66], stage07[68], stage06[71], stage05[72], stage04[88]}
   );
   gpc615_5 gpc615_5_107(
      {stage04[44], stage04[45], stage04[46], stage04[47], stage04[48]},
      {stage05[12]},
      {stage06[18], stage06[19], stage06[20], stage06[21], stage06[22], stage06[23]},
      {stage08[67], stage07[69], stage06[72], stage05[73], stage04[89]}
   );
   gpc615_5 gpc615_5_108(
      {stage04[49], stage04[50], stage04[51], stage04[52], stage04[53]},
      {stage05[13]},
      {stage06[24], stage06[25], stage06[26], stage06[27], stage06[28], stage06[29]},
      {stage08[68], stage07[70], stage06[73], stage05[74], stage04[90]}
   );
   gpc615_5 gpc615_5_109(
      {stage04[54], stage04[55], stage04[56], stage04[57], stage04[58]},
      {stage05[14]},
      {stage06[30], stage06[31], stage06[32], stage06[33], stage06[34], stage06[35]},
      {stage08[69], stage07[71], stage06[74], stage05[75], stage04[91]}
   );
   gpc615_5 gpc615_5_110(
      {stage04[59], stage04[60], stage04[61], stage04[62], stage04[63]},
      {stage05[15]},
      {stage06[36], stage06[37], stage06[38], stage06[39], stage06[40], stage06[41]},
      {stage08[70], stage07[72], stage06[75], stage05[76], stage04[92]}
   );
   gpc1_1 gpc1_1_111(
      {stage05[16]},
      {stage05[77]}
   );
   gpc1_1 gpc1_1_112(
      {stage05[17]},
      {stage05[78]}
   );
   gpc1_1 gpc1_1_113(
      {stage05[18]},
      {stage05[79]}
   );
   gpc1_1 gpc1_1_114(
      {stage05[19]},
      {stage05[80]}
   );
   gpc1_1 gpc1_1_115(
      {stage05[20]},
      {stage05[81]}
   );
   gpc1_1 gpc1_1_116(
      {stage05[21]},
      {stage05[82]}
   );
   gpc606_5 gpc606_5_117(
      {stage05[22], stage05[23], stage05[24], stage05[25], stage05[26], stage05[27]},
      {stage07[0], stage07[1], stage07[2], stage07[3], stage07[4], stage07[5]},
      {stage09[64], stage08[71], stage07[73], stage06[76], stage05[83]}
   );
   gpc606_5 gpc606_5_118(
      {stage05[28], stage05[29], stage05[30], stage05[31], stage05[32], stage05[33]},
      {stage07[6], stage07[7], stage07[8], stage07[9], stage07[10], stage07[11]},
      {stage09[65], stage08[72], stage07[74], stage06[77], stage05[84]}
   );
   gpc606_5 gpc606_5_119(
      {stage05[34], stage05[35], stage05[36], stage05[37], stage05[38], stage05[39]},
      {stage07[12], stage07[13], stage07[14], stage07[15], stage07[16], stage07[17]},
      {stage09[66], stage08[73], stage07[75], stage06[78], stage05[85]}
   );
   gpc606_5 gpc606_5_120(
      {stage05[40], stage05[41], stage05[42], stage05[43], stage05[44], stage05[45]},
      {stage07[18], stage07[19], stage07[20], stage07[21], stage07[22], stage07[23]},
      {stage09[67], stage08[74], stage07[76], stage06[79], stage05[86]}
   );
   gpc606_5 gpc606_5_121(
      {stage05[46], stage05[47], stage05[48], stage05[49], stage05[50], stage05[51]},
      {stage07[24], stage07[25], stage07[26], stage07[27], stage07[28], stage07[29]},
      {stage09[68], stage08[75], stage07[77], stage06[80], stage05[87]}
   );
   gpc606_5 gpc606_5_122(
      {stage05[52], stage05[53], stage05[54], stage05[55], stage05[56], stage05[57]},
      {stage07[30], stage07[31], stage07[32], stage07[33], stage07[34], stage07[35]},
      {stage09[69], stage08[76], stage07[78], stage06[81], stage05[88]}
   );
   gpc606_5 gpc606_5_123(
      {stage05[58], stage05[59], stage05[60], stage05[61], stage05[62], stage05[63]},
      {stage07[36], stage07[37], stage07[38], stage07[39], stage07[40], stage07[41]},
      {stage09[70], stage08[77], stage07[79], stage06[82], stage05[89]}
   );
   gpc1_1 gpc1_1_124(
      {stage06[42]},
      {stage06[83]}
   );
   gpc1_1 gpc1_1_125(
      {stage06[43]},
      {stage06[84]}
   );
   gpc1_1 gpc1_1_126(
      {stage06[44]},
      {stage06[85]}
   );
   gpc1_1 gpc1_1_127(
      {stage06[45]},
      {stage06[86]}
   );
   gpc606_5 gpc606_5_128(
      {stage06[46], stage06[47], stage06[48], stage06[49], stage06[50], stage06[51]},
      {stage08[0], stage08[1], stage08[2], stage08[3], stage08[4], stage08[5]},
      {stage10[64], stage09[71], stage08[78], stage07[80], stage06[87]}
   );
   gpc606_5 gpc606_5_129(
      {stage06[52], stage06[53], stage06[54], stage06[55], stage06[56], stage06[57]},
      {stage08[6], stage08[7], stage08[8], stage08[9], stage08[10], stage08[11]},
      {stage10[65], stage09[72], stage08[79], stage07[81], stage06[88]}
   );
   gpc606_5 gpc606_5_130(
      {stage06[58], stage06[59], stage06[60], stage06[61], stage06[62], stage06[63]},
      {stage08[12], stage08[13], stage08[14], stage08[15], stage08[16], stage08[17]},
      {stage10[66], stage09[73], stage08[80], stage07[82], stage06[89]}
   );
   gpc1_1 gpc1_1_131(
      {stage07[42]},
      {stage07[83]}
   );
   gpc1_1 gpc1_1_132(
      {stage07[43]},
      {stage07[84]}
   );
   gpc1_1 gpc1_1_133(
      {stage07[44]},
      {stage07[85]}
   );
   gpc1_1 gpc1_1_134(
      {stage07[45]},
      {stage07[86]}
   );
   gpc1_1 gpc1_1_135(
      {stage07[46]},
      {stage07[87]}
   );
   gpc1_1 gpc1_1_136(
      {stage07[47]},
      {stage07[88]}
   );
   gpc1_1 gpc1_1_137(
      {stage07[48]},
      {stage07[89]}
   );
   gpc1_1 gpc1_1_138(
      {stage07[49]},
      {stage07[90]}
   );
   gpc1_1 gpc1_1_139(
      {stage07[50]},
      {stage07[91]}
   );
   gpc1_1 gpc1_1_140(
      {stage07[51]},
      {stage07[92]}
   );
   gpc1_1 gpc1_1_141(
      {stage07[52]},
      {stage07[93]}
   );
   gpc1_1 gpc1_1_142(
      {stage07[53]},
      {stage07[94]}
   );
   gpc615_5 gpc615_5_143(
      {stage07[54], stage07[55], stage07[56], stage07[57], stage07[58]},
      {stage08[18]},
      {stage09[0], stage09[1], stage09[2], stage09[3], stage09[4], stage09[5]},
      {stage11[64], stage10[67], stage09[74], stage08[81], stage07[95]}
   );
   gpc615_5 gpc615_5_144(
      {stage07[59], stage07[60], stage07[61], stage07[62], stage07[63]},
      {stage08[19]},
      {stage09[6], stage09[7], stage09[8], stage09[9], stage09[10], stage09[11]},
      {stage11[65], stage10[68], stage09[75], stage08[82], stage07[96]}
   );
   gpc1_1 gpc1_1_145(
      {stage08[20]},
      {stage08[83]}
   );
   gpc1_1 gpc1_1_146(
      {stage08[21]},
      {stage08[84]}
   );
   gpc1_1 gpc1_1_147(
      {stage08[22]},
      {stage08[85]}
   );
   gpc1_1 gpc1_1_148(
      {stage08[23]},
      {stage08[86]}
   );
   gpc1_1 gpc1_1_149(
      {stage08[24]},
      {stage08[87]}
   );
   gpc1_1 gpc1_1_150(
      {stage08[25]},
      {stage08[88]}
   );
   gpc1_1 gpc1_1_151(
      {stage08[26]},
      {stage08[89]}
   );
   gpc1_1 gpc1_1_152(
      {stage08[27]},
      {stage08[90]}
   );
   gpc1_1 gpc1_1_153(
      {stage08[28]},
      {stage08[91]}
   );
   gpc1_1 gpc1_1_154(
      {stage08[29]},
      {stage08[92]}
   );
   gpc1_1 gpc1_1_155(
      {stage08[30]},
      {stage08[93]}
   );
   gpc1_1 gpc1_1_156(
      {stage08[31]},
      {stage08[94]}
   );
   gpc1_1 gpc1_1_157(
      {stage08[32]},
      {stage08[95]}
   );
   gpc1_1 gpc1_1_158(
      {stage08[33]},
      {stage08[96]}
   );
   gpc606_5 gpc606_5_159(
      {stage08[34], stage08[35], stage08[36], stage08[37], stage08[38], stage08[39]},
      {stage10[0], stage10[1], stage10[2], stage10[3], stage10[4], stage10[5]},
      {stage12[64], stage11[66], stage10[69], stage09[76], stage08[97]}
   );
   gpc606_5 gpc606_5_160(
      {stage08[40], stage08[41], stage08[42], stage08[43], stage08[44], stage08[45]},
      {stage10[6], stage10[7], stage10[8], stage10[9], stage10[10], stage10[11]},
      {stage12[65], stage11[67], stage10[70], stage09[77], stage08[98]}
   );
   gpc606_5 gpc606_5_161(
      {stage08[46], stage08[47], stage08[48], stage08[49], stage08[50], stage08[51]},
      {stage10[12], stage10[13], stage10[14], stage10[15], stage10[16], stage10[17]},
      {stage12[66], stage11[68], stage10[71], stage09[78], stage08[99]}
   );
   gpc606_5 gpc606_5_162(
      {stage08[52], stage08[53], stage08[54], stage08[55], stage08[56], stage08[57]},
      {stage10[18], stage10[19], stage10[20], stage10[21], stage10[22], stage10[23]},
      {stage12[67], stage11[69], stage10[72], stage09[79], stage08[100]}
   );
   gpc606_5 gpc606_5_163(
      {stage08[58], stage08[59], stage08[60], stage08[61], stage08[62], stage08[63]},
      {stage10[24], stage10[25], stage10[26], stage10[27], stage10[28], stage10[29]},
      {stage12[68], stage11[70], stage10[73], stage09[80], stage08[101]}
   );
   gpc1_1 gpc1_1_164(
      {stage09[12]},
      {stage09[81]}
   );
   gpc1_1 gpc1_1_165(
      {stage09[13]},
      {stage09[82]}
   );
   gpc1_1 gpc1_1_166(
      {stage09[14]},
      {stage09[83]}
   );
   gpc1_1 gpc1_1_167(
      {stage09[15]},
      {stage09[84]}
   );
   gpc1_1 gpc1_1_168(
      {stage09[16]},
      {stage09[85]}
   );
   gpc1_1 gpc1_1_169(
      {stage09[17]},
      {stage09[86]}
   );
   gpc1_1 gpc1_1_170(
      {stage09[18]},
      {stage09[87]}
   );
   gpc1_1 gpc1_1_171(
      {stage09[19]},
      {stage09[88]}
   );
   gpc1_1 gpc1_1_172(
      {stage09[20]},
      {stage09[89]}
   );
   gpc1_1 gpc1_1_173(
      {stage09[21]},
      {stage09[90]}
   );
   gpc1_1 gpc1_1_174(
      {stage09[22]},
      {stage09[91]}
   );
   gpc1_1 gpc1_1_175(
      {stage09[23]},
      {stage09[92]}
   );
   gpc1_1 gpc1_1_176(
      {stage09[24]},
      {stage09[93]}
   );
   gpc1_1 gpc1_1_177(
      {stage09[25]},
      {stage09[94]}
   );
   gpc1_1 gpc1_1_178(
      {stage09[26]},
      {stage09[95]}
   );
   gpc1_1 gpc1_1_179(
      {stage09[27]},
      {stage09[96]}
   );
   gpc1_1 gpc1_1_180(
      {stage09[28]},
      {stage09[97]}
   );
   gpc1_1 gpc1_1_181(
      {stage09[29]},
      {stage09[98]}
   );
   gpc1_1 gpc1_1_182(
      {stage09[30]},
      {stage09[99]}
   );
   gpc1_1 gpc1_1_183(
      {stage09[31]},
      {stage09[100]}
   );
   gpc1_1 gpc1_1_184(
      {stage09[32]},
      {stage09[101]}
   );
   gpc1_1 gpc1_1_185(
      {stage09[33]},
      {stage09[102]}
   );
   gpc1_1 gpc1_1_186(
      {stage09[34]},
      {stage09[103]}
   );
   gpc1_1 gpc1_1_187(
      {stage09[35]},
      {stage09[104]}
   );
   gpc1_1 gpc1_1_188(
      {stage09[36]},
      {stage09[105]}
   );
   gpc1_1 gpc1_1_189(
      {stage09[37]},
      {stage09[106]}
   );
   gpc1_1 gpc1_1_190(
      {stage09[38]},
      {stage09[107]}
   );
   gpc1_1 gpc1_1_191(
      {stage09[39]},
      {stage09[108]}
   );
   gpc1_1 gpc1_1_192(
      {stage09[40]},
      {stage09[109]}
   );
   gpc1_1 gpc1_1_193(
      {stage09[41]},
      {stage09[110]}
   );
   gpc1_1 gpc1_1_194(
      {stage09[42]},
      {stage09[111]}
   );
   gpc1_1 gpc1_1_195(
      {stage09[43]},
      {stage09[112]}
   );
   gpc1_1 gpc1_1_196(
      {stage09[44]},
      {stage09[113]}
   );
   gpc1_1 gpc1_1_197(
      {stage09[45]},
      {stage09[114]}
   );
   gpc1_1 gpc1_1_198(
      {stage09[46]},
      {stage09[115]}
   );
   gpc1_1 gpc1_1_199(
      {stage09[47]},
      {stage09[116]}
   );
   gpc1_1 gpc1_1_200(
      {stage09[48]},
      {stage09[117]}
   );
   gpc1_1 gpc1_1_201(
      {stage09[49]},
      {stage09[118]}
   );
   gpc1_1 gpc1_1_202(
      {stage09[50]},
      {stage09[119]}
   );
   gpc1_1 gpc1_1_203(
      {stage09[51]},
      {stage09[120]}
   );
   gpc606_5 gpc606_5_204(
      {stage09[52], stage09[53], stage09[54], stage09[55], stage09[56], stage09[57]},
      {stage11[0], stage11[1], stage11[2], stage11[3], stage11[4], stage11[5]},
      {stage13[64], stage12[69], stage11[71], stage10[74], stage09[121]}
   );
   gpc606_5 gpc606_5_205(
      {stage09[58], stage09[59], stage09[60], stage09[61], stage09[62], stage09[63]},
      {stage11[6], stage11[7], stage11[8], stage11[9], stage11[10], stage11[11]},
      {stage13[65], stage12[70], stage11[72], stage10[75], stage09[122]}
   );
   gpc1_1 gpc1_1_206(
      {stage10[30]},
      {stage10[76]}
   );
   gpc1_1 gpc1_1_207(
      {stage10[31]},
      {stage10[77]}
   );
   gpc1_1 gpc1_1_208(
      {stage10[32]},
      {stage10[78]}
   );
   gpc1_1 gpc1_1_209(
      {stage10[33]},
      {stage10[79]}
   );
   gpc1_1 gpc1_1_210(
      {stage10[34]},
      {stage10[80]}
   );
   gpc1_1 gpc1_1_211(
      {stage10[35]},
      {stage10[81]}
   );
   gpc1_1 gpc1_1_212(
      {stage10[36]},
      {stage10[82]}
   );
   gpc1_1 gpc1_1_213(
      {stage10[37]},
      {stage10[83]}
   );
   gpc1_1 gpc1_1_214(
      {stage10[38]},
      {stage10[84]}
   );
   gpc1_1 gpc1_1_215(
      {stage10[39]},
      {stage10[85]}
   );
   gpc1_1 gpc1_1_216(
      {stage10[40]},
      {stage10[86]}
   );
   gpc1_1 gpc1_1_217(
      {stage10[41]},
      {stage10[87]}
   );
   gpc1_1 gpc1_1_218(
      {stage10[42]},
      {stage10[88]}
   );
   gpc1_1 gpc1_1_219(
      {stage10[43]},
      {stage10[89]}
   );
   gpc1_1 gpc1_1_220(
      {stage10[44]},
      {stage10[90]}
   );
   gpc1_1 gpc1_1_221(
      {stage10[45]},
      {stage10[91]}
   );
   gpc1_1 gpc1_1_222(
      {stage10[46]},
      {stage10[92]}
   );
   gpc1_1 gpc1_1_223(
      {stage10[47]},
      {stage10[93]}
   );
   gpc1_1 gpc1_1_224(
      {stage10[48]},
      {stage10[94]}
   );
   gpc1_1 gpc1_1_225(
      {stage10[49]},
      {stage10[95]}
   );
   gpc1_1 gpc1_1_226(
      {stage10[50]},
      {stage10[96]}
   );
   gpc1_1 gpc1_1_227(
      {stage10[51]},
      {stage10[97]}
   );
   gpc1_1 gpc1_1_228(
      {stage10[52]},
      {stage10[98]}
   );
   gpc1_1 gpc1_1_229(
      {stage10[53]},
      {stage10[99]}
   );
   gpc1_1 gpc1_1_230(
      {stage10[54]},
      {stage10[100]}
   );
   gpc1_1 gpc1_1_231(
      {stage10[55]},
      {stage10[101]}
   );
   gpc1_1 gpc1_1_232(
      {stage10[56]},
      {stage10[102]}
   );
   gpc1_1 gpc1_1_233(
      {stage10[57]},
      {stage10[103]}
   );
   gpc1_1 gpc1_1_234(
      {stage10[58]},
      {stage10[104]}
   );
   gpc1_1 gpc1_1_235(
      {stage10[59]},
      {stage10[105]}
   );
   gpc1_1 gpc1_1_236(
      {stage10[60]},
      {stage10[106]}
   );
   gpc1_1 gpc1_1_237(
      {stage10[61]},
      {stage10[107]}
   );
   gpc1_1 gpc1_1_238(
      {stage10[62]},
      {stage10[108]}
   );
   gpc1_1 gpc1_1_239(
      {stage10[63]},
      {stage10[109]}
   );
   gpc1_1 gpc1_1_240(
      {stage11[12]},
      {stage11[73]}
   );
   gpc1_1 gpc1_1_241(
      {stage11[13]},
      {stage11[74]}
   );
   gpc1_1 gpc1_1_242(
      {stage11[14]},
      {stage11[75]}
   );
   gpc1_1 gpc1_1_243(
      {stage11[15]},
      {stage11[76]}
   );
   gpc1_1 gpc1_1_244(
      {stage11[16]},
      {stage11[77]}
   );
   gpc1_1 gpc1_1_245(
      {stage11[17]},
      {stage11[78]}
   );
   gpc1_1 gpc1_1_246(
      {stage11[18]},
      {stage11[79]}
   );
   gpc1_1 gpc1_1_247(
      {stage11[19]},
      {stage11[80]}
   );
   gpc1_1 gpc1_1_248(
      {stage11[20]},
      {stage11[81]}
   );
   gpc1_1 gpc1_1_249(
      {stage11[21]},
      {stage11[82]}
   );
   gpc1_1 gpc1_1_250(
      {stage11[22]},
      {stage11[83]}
   );
   gpc1_1 gpc1_1_251(
      {stage11[23]},
      {stage11[84]}
   );
   gpc615_5 gpc615_5_252(
      {stage11[24], stage11[25], stage11[26], stage11[27], stage11[28]},
      {stage12[0]},
      {stage13[0], stage13[1], stage13[2], stage13[3], stage13[4], stage13[5]},
      {stage15[64], stage14[64], stage13[66], stage12[71], stage11[85]}
   );
   gpc615_5 gpc615_5_253(
      {stage11[29], stage11[30], stage11[31], stage11[32], stage11[33]},
      {stage12[1]},
      {stage13[6], stage13[7], stage13[8], stage13[9], stage13[10], stage13[11]},
      {stage15[65], stage14[65], stage13[67], stage12[72], stage11[86]}
   );
   gpc615_5 gpc615_5_254(
      {stage11[34], stage11[35], stage11[36], stage11[37], stage11[38]},
      {stage12[2]},
      {stage13[12], stage13[13], stage13[14], stage13[15], stage13[16], stage13[17]},
      {stage15[66], stage14[66], stage13[68], stage12[73], stage11[87]}
   );
   gpc615_5 gpc615_5_255(
      {stage11[39], stage11[40], stage11[41], stage11[42], stage11[43]},
      {stage12[3]},
      {stage13[18], stage13[19], stage13[20], stage13[21], stage13[22], stage13[23]},
      {stage15[67], stage14[67], stage13[69], stage12[74], stage11[88]}
   );
   gpc615_5 gpc615_5_256(
      {stage11[44], stage11[45], stage11[46], stage11[47], stage11[48]},
      {stage12[4]},
      {stage13[24], stage13[25], stage13[26], stage13[27], stage13[28], stage13[29]},
      {stage15[68], stage14[68], stage13[70], stage12[75], stage11[89]}
   );
   gpc615_5 gpc615_5_257(
      {stage11[49], stage11[50], stage11[51], stage11[52], stage11[53]},
      {stage12[5]},
      {stage13[30], stage13[31], stage13[32], stage13[33], stage13[34], stage13[35]},
      {stage15[69], stage14[69], stage13[71], stage12[76], stage11[90]}
   );
   gpc615_5 gpc615_5_258(
      {stage11[54], stage11[55], stage11[56], stage11[57], stage11[58]},
      {stage12[6]},
      {stage13[36], stage13[37], stage13[38], stage13[39], stage13[40], stage13[41]},
      {stage15[70], stage14[70], stage13[72], stage12[77], stage11[91]}
   );
   gpc615_5 gpc615_5_259(
      {stage11[59], stage11[60], stage11[61], stage11[62], stage11[63]},
      {stage12[7]},
      {stage13[42], stage13[43], stage13[44], stage13[45], stage13[46], stage13[47]},
      {stage15[71], stage14[71], stage13[73], stage12[78], stage11[92]}
   );
   gpc1_1 gpc1_1_260(
      {stage12[8]},
      {stage12[79]}
   );
   gpc1_1 gpc1_1_261(
      {stage12[9]},
      {stage12[80]}
   );
   gpc1_1 gpc1_1_262(
      {stage12[10]},
      {stage12[81]}
   );
   gpc1_1 gpc1_1_263(
      {stage12[11]},
      {stage12[82]}
   );
   gpc1_1 gpc1_1_264(
      {stage12[12]},
      {stage12[83]}
   );
   gpc1_1 gpc1_1_265(
      {stage12[13]},
      {stage12[84]}
   );
   gpc1_1 gpc1_1_266(
      {stage12[14]},
      {stage12[85]}
   );
   gpc1_1 gpc1_1_267(
      {stage12[15]},
      {stage12[86]}
   );
   gpc1_1 gpc1_1_268(
      {stage12[16]},
      {stage12[87]}
   );
   gpc1_1 gpc1_1_269(
      {stage12[17]},
      {stage12[88]}
   );
   gpc1_1 gpc1_1_270(
      {stage12[18]},
      {stage12[89]}
   );
   gpc1_1 gpc1_1_271(
      {stage12[19]},
      {stage12[90]}
   );
   gpc1_1 gpc1_1_272(
      {stage12[20]},
      {stage12[91]}
   );
   gpc1_1 gpc1_1_273(
      {stage12[21]},
      {stage12[92]}
   );
   gpc1_1 gpc1_1_274(
      {stage12[22]},
      {stage12[93]}
   );
   gpc1_1 gpc1_1_275(
      {stage12[23]},
      {stage12[94]}
   );
   gpc1_1 gpc1_1_276(
      {stage12[24]},
      {stage12[95]}
   );
   gpc1_1 gpc1_1_277(
      {stage12[25]},
      {stage12[96]}
   );
   gpc1_1 gpc1_1_278(
      {stage12[26]},
      {stage12[97]}
   );
   gpc1_1 gpc1_1_279(
      {stage12[27]},
      {stage12[98]}
   );
   gpc1_1 gpc1_1_280(
      {stage12[28]},
      {stage12[99]}
   );
   gpc1_1 gpc1_1_281(
      {stage12[29]},
      {stage12[100]}
   );
   gpc1_1 gpc1_1_282(
      {stage12[30]},
      {stage12[101]}
   );
   gpc1_1 gpc1_1_283(
      {stage12[31]},
      {stage12[102]}
   );
   gpc1_1 gpc1_1_284(
      {stage12[32]},
      {stage12[103]}
   );
   gpc1_1 gpc1_1_285(
      {stage12[33]},
      {stage12[104]}
   );
   gpc606_5 gpc606_5_286(
      {stage12[34], stage12[35], stage12[36], stage12[37], stage12[38], stage12[39]},
      {stage14[0], stage14[1], stage14[2], stage14[3], stage14[4], stage14[5]},
      {stage16[64], stage15[72], stage14[72], stage13[74], stage12[105]}
   );
   gpc606_5 gpc606_5_287(
      {stage12[40], stage12[41], stage12[42], stage12[43], stage12[44], stage12[45]},
      {stage14[6], stage14[7], stage14[8], stage14[9], stage14[10], stage14[11]},
      {stage16[65], stage15[73], stage14[73], stage13[75], stage12[106]}
   );
   gpc606_5 gpc606_5_288(
      {stage12[46], stage12[47], stage12[48], stage12[49], stage12[50], stage12[51]},
      {stage14[12], stage14[13], stage14[14], stage14[15], stage14[16], stage14[17]},
      {stage16[66], stage15[74], stage14[74], stage13[76], stage12[107]}
   );
   gpc606_5 gpc606_5_289(
      {stage12[52], stage12[53], stage12[54], stage12[55], stage12[56], stage12[57]},
      {stage14[18], stage14[19], stage14[20], stage14[21], stage14[22], stage14[23]},
      {stage16[67], stage15[75], stage14[75], stage13[77], stage12[108]}
   );
   gpc606_5 gpc606_5_290(
      {stage12[58], stage12[59], stage12[60], stage12[61], stage12[62], stage12[63]},
      {stage14[24], stage14[25], stage14[26], stage14[27], stage14[28], stage14[29]},
      {stage16[68], stage15[76], stage14[76], stage13[78], stage12[109]}
   );
   gpc1_1 gpc1_1_291(
      {stage13[48]},
      {stage13[79]}
   );
   gpc1_1 gpc1_1_292(
      {stage13[49]},
      {stage13[80]}
   );
   gpc1_1 gpc1_1_293(
      {stage13[50]},
      {stage13[81]}
   );
   gpc1_1 gpc1_1_294(
      {stage13[51]},
      {stage13[82]}
   );
   gpc1_1 gpc1_1_295(
      {stage13[52]},
      {stage13[83]}
   );
   gpc1_1 gpc1_1_296(
      {stage13[53]},
      {stage13[84]}
   );
   gpc1_1 gpc1_1_297(
      {stage13[54]},
      {stage13[85]}
   );
   gpc1_1 gpc1_1_298(
      {stage13[55]},
      {stage13[86]}
   );
   gpc1_1 gpc1_1_299(
      {stage13[56]},
      {stage13[87]}
   );
   gpc1_1 gpc1_1_300(
      {stage13[57]},
      {stage13[88]}
   );
   gpc606_5 gpc606_5_301(
      {stage13[58], stage13[59], stage13[60], stage13[61], stage13[62], stage13[63]},
      {stage15[0], stage15[1], stage15[2], stage15[3], stage15[4], stage15[5]},
      {stage17[64], stage16[69], stage15[77], stage14[77], stage13[89]}
   );
   gpc1_1 gpc1_1_302(
      {stage14[30]},
      {stage14[78]}
   );
   gpc1_1 gpc1_1_303(
      {stage14[31]},
      {stage14[79]}
   );
   gpc1_1 gpc1_1_304(
      {stage14[32]},
      {stage14[80]}
   );
   gpc1_1 gpc1_1_305(
      {stage14[33]},
      {stage14[81]}
   );
   gpc1_1 gpc1_1_306(
      {stage14[34]},
      {stage14[82]}
   );
   gpc1_1 gpc1_1_307(
      {stage14[35]},
      {stage14[83]}
   );
   gpc1_1 gpc1_1_308(
      {stage14[36]},
      {stage14[84]}
   );
   gpc1_1 gpc1_1_309(
      {stage14[37]},
      {stage14[85]}
   );
   gpc1_1 gpc1_1_310(
      {stage14[38]},
      {stage14[86]}
   );
   gpc1_1 gpc1_1_311(
      {stage14[39]},
      {stage14[87]}
   );
   gpc1_1 gpc1_1_312(
      {stage14[40]},
      {stage14[88]}
   );
   gpc1_1 gpc1_1_313(
      {stage14[41]},
      {stage14[89]}
   );
   gpc1_1 gpc1_1_314(
      {stage14[42]},
      {stage14[90]}
   );
   gpc7_3 gpc7_3_315(
      {stage14[43], stage14[44], stage14[45], stage14[46], stage14[47], stage14[48], stage14[49]},
      {stage16[70], stage15[78], stage14[91]}
   );
   gpc7_3 gpc7_3_316(
      {stage14[50], stage14[51], stage14[52], stage14[53], stage14[54], stage14[55], stage14[56]},
      {stage16[71], stage15[79], stage14[92]}
   );
   gpc7_3 gpc7_3_317(
      {stage14[57], stage14[58], stage14[59], stage14[60], stage14[61], stage14[62], stage14[63]},
      {stage16[72], stage15[80], stage14[93]}
   );
   gpc1_1 gpc1_1_318(
      {stage15[6]},
      {stage15[81]}
   );
   gpc1_1 gpc1_1_319(
      {stage15[7]},
      {stage15[82]}
   );
   gpc1_1 gpc1_1_320(
      {stage15[8]},
      {stage15[83]}
   );
   gpc1_1 gpc1_1_321(
      {stage15[9]},
      {stage15[84]}
   );
   gpc1_1 gpc1_1_322(
      {stage15[10]},
      {stage15[85]}
   );
   gpc1_1 gpc1_1_323(
      {stage15[11]},
      {stage15[86]}
   );
   gpc1_1 gpc1_1_324(
      {stage15[12]},
      {stage15[87]}
   );
   gpc1_1 gpc1_1_325(
      {stage15[13]},
      {stage15[88]}
   );
   gpc1_1 gpc1_1_326(
      {stage15[14]},
      {stage15[89]}
   );
   gpc1_1 gpc1_1_327(
      {stage15[15]},
      {stage15[90]}
   );
   gpc1_1 gpc1_1_328(
      {stage15[16]},
      {stage15[91]}
   );
   gpc1_1 gpc1_1_329(
      {stage15[17]},
      {stage15[92]}
   );
   gpc1_1 gpc1_1_330(
      {stage15[18]},
      {stage15[93]}
   );
   gpc1_1 gpc1_1_331(
      {stage15[19]},
      {stage15[94]}
   );
   gpc1_1 gpc1_1_332(
      {stage15[20]},
      {stage15[95]}
   );
   gpc1_1 gpc1_1_333(
      {stage15[21]},
      {stage15[96]}
   );
   gpc1_1 gpc1_1_334(
      {stage15[22]},
      {stage15[97]}
   );
   gpc1_1 gpc1_1_335(
      {stage15[23]},
      {stage15[98]}
   );
   gpc1_1 gpc1_1_336(
      {stage15[24]},
      {stage15[99]}
   );
   gpc1_1 gpc1_1_337(
      {stage15[25]},
      {stage15[100]}
   );
   gpc1_1 gpc1_1_338(
      {stage15[26]},
      {stage15[101]}
   );
   gpc1_1 gpc1_1_339(
      {stage15[27]},
      {stage15[102]}
   );
   gpc1_1 gpc1_1_340(
      {stage15[28]},
      {stage15[103]}
   );
   gpc1_1 gpc1_1_341(
      {stage15[29]},
      {stage15[104]}
   );
   gpc1_1 gpc1_1_342(
      {stage15[30]},
      {stage15[105]}
   );
   gpc1_1 gpc1_1_343(
      {stage15[31]},
      {stage15[106]}
   );
   gpc1_1 gpc1_1_344(
      {stage15[32]},
      {stage15[107]}
   );
   gpc1_1 gpc1_1_345(
      {stage15[33]},
      {stage15[108]}
   );
   gpc1_1 gpc1_1_346(
      {stage15[34]},
      {stage15[109]}
   );
   gpc1_1 gpc1_1_347(
      {stage15[35]},
      {stage15[110]}
   );
   gpc1_1 gpc1_1_348(
      {stage15[36]},
      {stage15[111]}
   );
   gpc1_1 gpc1_1_349(
      {stage15[37]},
      {stage15[112]}
   );
   gpc1_1 gpc1_1_350(
      {stage15[38]},
      {stage15[113]}
   );
   gpc1_1 gpc1_1_351(
      {stage15[39]},
      {stage15[114]}
   );
   gpc1_1 gpc1_1_352(
      {stage15[40]},
      {stage15[115]}
   );
   gpc1_1 gpc1_1_353(
      {stage15[41]},
      {stage15[116]}
   );
   gpc1_1 gpc1_1_354(
      {stage15[42]},
      {stage15[117]}
   );
   gpc1_1 gpc1_1_355(
      {stage15[43]},
      {stage15[118]}
   );
   gpc1_1 gpc1_1_356(
      {stage15[44]},
      {stage15[119]}
   );
   gpc1_1 gpc1_1_357(
      {stage15[45]},
      {stage15[120]}
   );
   gpc606_5 gpc606_5_358(
      {stage15[46], stage15[47], stage15[48], stage15[49], stage15[50], stage15[51]},
      {stage17[0], stage17[1], stage17[2], stage17[3], stage17[4], stage17[5]},
      {stage19[64], stage18[64], stage17[65], stage16[73], stage15[121]}
   );
   gpc606_5 gpc606_5_359(
      {stage15[52], stage15[53], stage15[54], stage15[55], stage15[56], stage15[57]},
      {stage17[6], stage17[7], stage17[8], stage17[9], stage17[10], stage17[11]},
      {stage19[65], stage18[65], stage17[66], stage16[74], stage15[122]}
   );
   gpc606_5 gpc606_5_360(
      {stage15[58], stage15[59], stage15[60], stage15[61], stage15[62], stage15[63]},
      {stage17[12], stage17[13], stage17[14], stage17[15], stage17[16], stage17[17]},
      {stage19[66], stage18[66], stage17[67], stage16[75], stage15[123]}
   );
   gpc1_1 gpc1_1_361(
      {stage16[0]},
      {stage16[76]}
   );
   gpc1_1 gpc1_1_362(
      {stage16[1]},
      {stage16[77]}
   );
   gpc1_1 gpc1_1_363(
      {stage16[2]},
      {stage16[78]}
   );
   gpc1_1 gpc1_1_364(
      {stage16[3]},
      {stage16[79]}
   );
   gpc606_5 gpc606_5_365(
      {stage16[4], stage16[5], stage16[6], stage16[7], stage16[8], stage16[9]},
      {stage18[0], stage18[1], stage18[2], stage18[3], stage18[4], stage18[5]},
      {stage20[64], stage19[67], stage18[67], stage17[68], stage16[80]}
   );
   gpc606_5 gpc606_5_366(
      {stage16[10], stage16[11], stage16[12], stage16[13], stage16[14], stage16[15]},
      {stage18[6], stage18[7], stage18[8], stage18[9], stage18[10], stage18[11]},
      {stage20[65], stage19[68], stage18[68], stage17[69], stage16[81]}
   );
   gpc606_5 gpc606_5_367(
      {stage16[16], stage16[17], stage16[18], stage16[19], stage16[20], stage16[21]},
      {stage18[12], stage18[13], stage18[14], stage18[15], stage18[16], stage18[17]},
      {stage20[66], stage19[69], stage18[69], stage17[70], stage16[82]}
   );
   gpc606_5 gpc606_5_368(
      {stage16[22], stage16[23], stage16[24], stage16[25], stage16[26], stage16[27]},
      {stage18[18], stage18[19], stage18[20], stage18[21], stage18[22], stage18[23]},
      {stage20[67], stage19[70], stage18[70], stage17[71], stage16[83]}
   );
   gpc606_5 gpc606_5_369(
      {stage16[28], stage16[29], stage16[30], stage16[31], stage16[32], stage16[33]},
      {stage18[24], stage18[25], stage18[26], stage18[27], stage18[28], stage18[29]},
      {stage20[68], stage19[71], stage18[71], stage17[72], stage16[84]}
   );
   gpc606_5 gpc606_5_370(
      {stage16[34], stage16[35], stage16[36], stage16[37], stage16[38], stage16[39]},
      {stage18[30], stage18[31], stage18[32], stage18[33], stage18[34], stage18[35]},
      {stage20[69], stage19[72], stage18[72], stage17[73], stage16[85]}
   );
   gpc606_5 gpc606_5_371(
      {stage16[40], stage16[41], stage16[42], stage16[43], stage16[44], stage16[45]},
      {stage18[36], stage18[37], stage18[38], stage18[39], stage18[40], stage18[41]},
      {stage20[70], stage19[73], stage18[73], stage17[74], stage16[86]}
   );
   gpc606_5 gpc606_5_372(
      {stage16[46], stage16[47], stage16[48], stage16[49], stage16[50], stage16[51]},
      {stage18[42], stage18[43], stage18[44], stage18[45], stage18[46], stage18[47]},
      {stage20[71], stage19[74], stage18[74], stage17[75], stage16[87]}
   );
   gpc606_5 gpc606_5_373(
      {stage16[52], stage16[53], stage16[54], stage16[55], stage16[56], stage16[57]},
      {stage18[48], stage18[49], stage18[50], stage18[51], stage18[52], stage18[53]},
      {stage20[72], stage19[75], stage18[75], stage17[76], stage16[88]}
   );
   gpc606_5 gpc606_5_374(
      {stage16[58], stage16[59], stage16[60], stage16[61], stage16[62], stage16[63]},
      {stage18[54], stage18[55], stage18[56], stage18[57], stage18[58], stage18[59]},
      {stage20[73], stage19[76], stage18[76], stage17[77], stage16[89]}
   );
   gpc1_1 gpc1_1_375(
      {stage17[18]},
      {stage17[78]}
   );
   gpc1_1 gpc1_1_376(
      {stage17[19]},
      {stage17[79]}
   );
   gpc1_1 gpc1_1_377(
      {stage17[20]},
      {stage17[80]}
   );
   gpc1_1 gpc1_1_378(
      {stage17[21]},
      {stage17[81]}
   );
   gpc1_1 gpc1_1_379(
      {stage17[22]},
      {stage17[82]}
   );
   gpc1_1 gpc1_1_380(
      {stage17[23]},
      {stage17[83]}
   );
   gpc1_1 gpc1_1_381(
      {stage17[24]},
      {stage17[84]}
   );
   gpc1_1 gpc1_1_382(
      {stage17[25]},
      {stage17[85]}
   );
   gpc1_1 gpc1_1_383(
      {stage17[26]},
      {stage17[86]}
   );
   gpc1_1 gpc1_1_384(
      {stage17[27]},
      {stage17[87]}
   );
   gpc1_1 gpc1_1_385(
      {stage17[28]},
      {stage17[88]}
   );
   gpc1_1 gpc1_1_386(
      {stage17[29]},
      {stage17[89]}
   );
   gpc1_1 gpc1_1_387(
      {stage17[30]},
      {stage17[90]}
   );
   gpc1_1 gpc1_1_388(
      {stage17[31]},
      {stage17[91]}
   );
   gpc1_1 gpc1_1_389(
      {stage17[32]},
      {stage17[92]}
   );
   gpc1_1 gpc1_1_390(
      {stage17[33]},
      {stage17[93]}
   );
   gpc1_1 gpc1_1_391(
      {stage17[34]},
      {stage17[94]}
   );
   gpc1_1 gpc1_1_392(
      {stage17[35]},
      {stage17[95]}
   );
   gpc1_1 gpc1_1_393(
      {stage17[36]},
      {stage17[96]}
   );
   gpc1_1 gpc1_1_394(
      {stage17[37]},
      {stage17[97]}
   );
   gpc1_1 gpc1_1_395(
      {stage17[38]},
      {stage17[98]}
   );
   gpc1_1 gpc1_1_396(
      {stage17[39]},
      {stage17[99]}
   );
   gpc606_5 gpc606_5_397(
      {stage17[40], stage17[41], stage17[42], stage17[43], stage17[44], stage17[45]},
      {stage19[0], stage19[1], stage19[2], stage19[3], stage19[4], stage19[5]},
      {stage21[64], stage20[74], stage19[77], stage18[77], stage17[100]}
   );
   gpc606_5 gpc606_5_398(
      {stage17[46], stage17[47], stage17[48], stage17[49], stage17[50], stage17[51]},
      {stage19[6], stage19[7], stage19[8], stage19[9], stage19[10], stage19[11]},
      {stage21[65], stage20[75], stage19[78], stage18[78], stage17[101]}
   );
   gpc606_5 gpc606_5_399(
      {stage17[52], stage17[53], stage17[54], stage17[55], stage17[56], stage17[57]},
      {stage19[12], stage19[13], stage19[14], stage19[15], stage19[16], stage19[17]},
      {stage21[66], stage20[76], stage19[79], stage18[79], stage17[102]}
   );
   gpc1406_5 gpc1406_5_400(
      {stage17[58], stage17[59], stage17[60], stage17[61], stage17[62], stage17[63]},
      {stage19[18], stage19[19], stage19[20], stage19[21]},
      {stage20[0]},
      {stage21[67], stage20[77], stage19[80], stage18[80], stage17[103]}
   );
   gpc1_1 gpc1_1_401(
      {stage18[60]},
      {stage18[81]}
   );
   gpc1_1 gpc1_1_402(
      {stage18[61]},
      {stage18[82]}
   );
   gpc1_1 gpc1_1_403(
      {stage18[62]},
      {stage18[83]}
   );
   gpc1_1 gpc1_1_404(
      {stage18[63]},
      {stage18[84]}
   );
   gpc1_1 gpc1_1_405(
      {stage19[22]},
      {stage19[81]}
   );
   gpc1_1 gpc1_1_406(
      {stage19[23]},
      {stage19[82]}
   );
   gpc1_1 gpc1_1_407(
      {stage19[24]},
      {stage19[83]}
   );
   gpc1_1 gpc1_1_408(
      {stage19[25]},
      {stage19[84]}
   );
   gpc1_1 gpc1_1_409(
      {stage19[26]},
      {stage19[85]}
   );
   gpc1_1 gpc1_1_410(
      {stage19[27]},
      {stage19[86]}
   );
   gpc1_1 gpc1_1_411(
      {stage19[28]},
      {stage19[87]}
   );
   gpc1_1 gpc1_1_412(
      {stage19[29]},
      {stage19[88]}
   );
   gpc1_1 gpc1_1_413(
      {stage19[30]},
      {stage19[89]}
   );
   gpc1_1 gpc1_1_414(
      {stage19[31]},
      {stage19[90]}
   );
   gpc1_1 gpc1_1_415(
      {stage19[32]},
      {stage19[91]}
   );
   gpc1_1 gpc1_1_416(
      {stage19[33]},
      {stage19[92]}
   );
   gpc1_1 gpc1_1_417(
      {stage19[34]},
      {stage19[93]}
   );
   gpc606_5 gpc606_5_418(
      {stage19[35], stage19[36], stage19[37], stage19[38], stage19[39], stage19[40]},
      {stage21[0], stage21[1], stage21[2], stage21[3], stage21[4], stage21[5]},
      {stage23[64], stage22[64], stage21[68], stage20[78], stage19[94]}
   );
   gpc606_5 gpc606_5_419(
      {stage19[41], stage19[42], stage19[43], stage19[44], stage19[45], stage19[46]},
      {stage21[6], stage21[7], stage21[8], stage21[9], stage21[10], stage21[11]},
      {stage23[65], stage22[65], stage21[69], stage20[79], stage19[95]}
   );
   gpc606_5 gpc606_5_420(
      {stage19[47], stage19[48], stage19[49], stage19[50], stage19[51], stage19[52]},
      {stage21[12], stage21[13], stage21[14], stage21[15], stage21[16], stage21[17]},
      {stage23[66], stage22[66], stage21[70], stage20[80], stage19[96]}
   );
   gpc606_5 gpc606_5_421(
      {stage19[53], stage19[54], stage19[55], stage19[56], stage19[57], stage19[58]},
      {stage21[18], stage21[19], stage21[20], stage21[21], stage21[22], stage21[23]},
      {stage23[67], stage22[67], stage21[71], stage20[81], stage19[97]}
   );
   gpc215_4 gpc215_4_422(
      {stage19[59], stage19[60], stage19[61], stage19[62], stage19[63]},
      {stage20[1]},
      {stage21[24], stage21[25]},
      {stage22[68], stage21[72], stage20[82], stage19[98]}
   );
   gpc1_1 gpc1_1_423(
      {stage20[2]},
      {stage20[83]}
   );
   gpc1_1 gpc1_1_424(
      {stage20[3]},
      {stage20[84]}
   );
   gpc1_1 gpc1_1_425(
      {stage20[4]},
      {stage20[85]}
   );
   gpc1_1 gpc1_1_426(
      {stage20[5]},
      {stage20[86]}
   );
   gpc1_1 gpc1_1_427(
      {stage20[6]},
      {stage20[87]}
   );
   gpc1_1 gpc1_1_428(
      {stage20[7]},
      {stage20[88]}
   );
   gpc1_1 gpc1_1_429(
      {stage20[8]},
      {stage20[89]}
   );
   gpc1_1 gpc1_1_430(
      {stage20[9]},
      {stage20[90]}
   );
   gpc1_1 gpc1_1_431(
      {stage20[10]},
      {stage20[91]}
   );
   gpc1_1 gpc1_1_432(
      {stage20[11]},
      {stage20[92]}
   );
   gpc1_1 gpc1_1_433(
      {stage20[12]},
      {stage20[93]}
   );
   gpc1_1 gpc1_1_434(
      {stage20[13]},
      {stage20[94]}
   );
   gpc1_1 gpc1_1_435(
      {stage20[14]},
      {stage20[95]}
   );
   gpc1_1 gpc1_1_436(
      {stage20[15]},
      {stage20[96]}
   );
   gpc1_1 gpc1_1_437(
      {stage20[16]},
      {stage20[97]}
   );
   gpc606_5 gpc606_5_438(
      {stage20[17], stage20[18], stage20[19], stage20[20], stage20[21], stage20[22]},
      {stage22[0], stage22[1], stage22[2], stage22[3], stage22[4], stage22[5]},
      {stage24[64], stage23[68], stage22[69], stage21[73], stage20[98]}
   );
   gpc606_5 gpc606_5_439(
      {stage20[23], stage20[24], stage20[25], stage20[26], stage20[27], stage20[28]},
      {stage22[6], stage22[7], stage22[8], stage22[9], stage22[10], stage22[11]},
      {stage24[65], stage23[69], stage22[70], stage21[74], stage20[99]}
   );
   gpc606_5 gpc606_5_440(
      {stage20[29], stage20[30], stage20[31], stage20[32], stage20[33], stage20[34]},
      {stage22[12], stage22[13], stage22[14], stage22[15], stage22[16], stage22[17]},
      {stage24[66], stage23[70], stage22[71], stage21[75], stage20[100]}
   );
   gpc606_5 gpc606_5_441(
      {stage20[35], stage20[36], stage20[37], stage20[38], stage20[39], stage20[40]},
      {stage22[18], stage22[19], stage22[20], stage22[21], stage22[22], stage22[23]},
      {stage24[67], stage23[71], stage22[72], stage21[76], stage20[101]}
   );
   gpc606_5 gpc606_5_442(
      {stage20[41], stage20[42], stage20[43], stage20[44], stage20[45], stage20[46]},
      {stage22[24], stage22[25], stage22[26], stage22[27], stage22[28], stage22[29]},
      {stage24[68], stage23[72], stage22[73], stage21[77], stage20[102]}
   );
   gpc606_5 gpc606_5_443(
      {stage20[47], stage20[48], stage20[49], stage20[50], stage20[51], stage20[52]},
      {stage22[30], stage22[31], stage22[32], stage22[33], stage22[34], stage22[35]},
      {stage24[69], stage23[73], stage22[74], stage21[78], stage20[103]}
   );
   gpc606_5 gpc606_5_444(
      {stage20[53], stage20[54], stage20[55], stage20[56], stage20[57], stage20[58]},
      {stage22[36], stage22[37], stage22[38], stage22[39], stage22[40], stage22[41]},
      {stage24[70], stage23[74], stage22[75], stage21[79], stage20[104]}
   );
   gpc2135_5 gpc2135_5_445(
      {stage20[59], stage20[60], stage20[61], stage20[62], stage20[63]},
      {stage21[26], stage21[27], stage21[28]},
      {stage22[42]},
      {stage23[0], stage23[1]},
      {stage24[71], stage23[75], stage22[76], stage21[80], stage20[105]}
   );
   gpc1_1 gpc1_1_446(
      {stage21[29]},
      {stage21[81]}
   );
   gpc1_1 gpc1_1_447(
      {stage21[30]},
      {stage21[82]}
   );
   gpc1_1 gpc1_1_448(
      {stage21[31]},
      {stage21[83]}
   );
   gpc1_1 gpc1_1_449(
      {stage21[32]},
      {stage21[84]}
   );
   gpc1_1 gpc1_1_450(
      {stage21[33]},
      {stage21[85]}
   );
   gpc606_5 gpc606_5_451(
      {stage21[34], stage21[35], stage21[36], stage21[37], stage21[38], stage21[39]},
      {stage23[2], stage23[3], stage23[4], stage23[5], stage23[6], stage23[7]},
      {stage25[64], stage24[72], stage23[76], stage22[77], stage21[86]}
   );
   gpc606_5 gpc606_5_452(
      {stage21[40], stage21[41], stage21[42], stage21[43], stage21[44], stage21[45]},
      {stage23[8], stage23[9], stage23[10], stage23[11], stage23[12], stage23[13]},
      {stage25[65], stage24[73], stage23[77], stage22[78], stage21[87]}
   );
   gpc606_5 gpc606_5_453(
      {stage21[46], stage21[47], stage21[48], stage21[49], stage21[50], stage21[51]},
      {stage23[14], stage23[15], stage23[16], stage23[17], stage23[18], stage23[19]},
      {stage25[66], stage24[74], stage23[78], stage22[79], stage21[88]}
   );
   gpc606_5 gpc606_5_454(
      {stage21[52], stage21[53], stage21[54], stage21[55], stage21[56], stage21[57]},
      {stage23[20], stage23[21], stage23[22], stage23[23], stage23[24], stage23[25]},
      {stage25[67], stage24[75], stage23[79], stage22[80], stage21[89]}
   );
   gpc606_5 gpc606_5_455(
      {stage21[58], stage21[59], stage21[60], stage21[61], stage21[62], stage21[63]},
      {stage23[26], stage23[27], stage23[28], stage23[29], stage23[30], stage23[31]},
      {stage25[68], stage24[76], stage23[80], stage22[81], stage21[90]}
   );
   gpc1_1 gpc1_1_456(
      {stage22[43]},
      {stage22[82]}
   );
   gpc1_1 gpc1_1_457(
      {stage22[44]},
      {stage22[83]}
   );
   gpc1_1 gpc1_1_458(
      {stage22[45]},
      {stage22[84]}
   );
   gpc1_1 gpc1_1_459(
      {stage22[46]},
      {stage22[85]}
   );
   gpc1_1 gpc1_1_460(
      {stage22[47]},
      {stage22[86]}
   );
   gpc1_1 gpc1_1_461(
      {stage22[48]},
      {stage22[87]}
   );
   gpc1_1 gpc1_1_462(
      {stage22[49]},
      {stage22[88]}
   );
   gpc1_1 gpc1_1_463(
      {stage22[50]},
      {stage22[89]}
   );
   gpc1_1 gpc1_1_464(
      {stage22[51]},
      {stage22[90]}
   );
   gpc1_1 gpc1_1_465(
      {stage22[52]},
      {stage22[91]}
   );
   gpc1_1 gpc1_1_466(
      {stage22[53]},
      {stage22[92]}
   );
   gpc1_1 gpc1_1_467(
      {stage22[54]},
      {stage22[93]}
   );
   gpc1_1 gpc1_1_468(
      {stage22[55]},
      {stage22[94]}
   );
   gpc1_1 gpc1_1_469(
      {stage22[56]},
      {stage22[95]}
   );
   gpc1_1 gpc1_1_470(
      {stage22[57]},
      {stage22[96]}
   );
   gpc1_1 gpc1_1_471(
      {stage22[58]},
      {stage22[97]}
   );
   gpc615_5 gpc615_5_472(
      {stage22[59], stage22[60], stage22[61], stage22[62], stage22[63]},
      {stage23[32]},
      {stage24[0], stage24[1], stage24[2], stage24[3], stage24[4], stage24[5]},
      {stage26[64], stage25[69], stage24[77], stage23[81], stage22[98]}
   );
   gpc1_1 gpc1_1_473(
      {stage23[33]},
      {stage23[82]}
   );
   gpc1_1 gpc1_1_474(
      {stage23[34]},
      {stage23[83]}
   );
   gpc1_1 gpc1_1_475(
      {stage23[35]},
      {stage23[84]}
   );
   gpc1_1 gpc1_1_476(
      {stage23[36]},
      {stage23[85]}
   );
   gpc1_1 gpc1_1_477(
      {stage23[37]},
      {stage23[86]}
   );
   gpc1_1 gpc1_1_478(
      {stage23[38]},
      {stage23[87]}
   );
   gpc1_1 gpc1_1_479(
      {stage23[39]},
      {stage23[88]}
   );
   gpc1_1 gpc1_1_480(
      {stage23[40]},
      {stage23[89]}
   );
   gpc1_1 gpc1_1_481(
      {stage23[41]},
      {stage23[90]}
   );
   gpc7_3 gpc7_3_482(
      {stage23[42], stage23[43], stage23[44], stage23[45], stage23[46], stage23[47], stage23[48]},
      {stage25[70], stage24[78], stage23[91]}
   );
   gpc615_5 gpc615_5_483(
      {stage23[49], stage23[50], stage23[51], stage23[52], stage23[53]},
      {stage24[6]},
      {stage25[0], stage25[1], stage25[2], stage25[3], stage25[4], stage25[5]},
      {stage27[64], stage26[65], stage25[71], stage24[79], stage23[92]}
   );
   gpc615_5 gpc615_5_484(
      {stage23[54], stage23[55], stage23[56], stage23[57], stage23[58]},
      {stage24[7]},
      {stage25[6], stage25[7], stage25[8], stage25[9], stage25[10], stage25[11]},
      {stage27[65], stage26[66], stage25[72], stage24[80], stage23[93]}
   );
   gpc615_5 gpc615_5_485(
      {stage23[59], stage23[60], stage23[61], stage23[62], stage23[63]},
      {stage24[8]},
      {stage25[12], stage25[13], stage25[14], stage25[15], stage25[16], stage25[17]},
      {stage27[66], stage26[67], stage25[73], stage24[81], stage23[94]}
   );
   gpc1_1 gpc1_1_486(
      {stage24[9]},
      {stage24[82]}
   );
   gpc1_1 gpc1_1_487(
      {stage24[10]},
      {stage24[83]}
   );
   gpc1_1 gpc1_1_488(
      {stage24[11]},
      {stage24[84]}
   );
   gpc1_1 gpc1_1_489(
      {stage24[12]},
      {stage24[85]}
   );
   gpc1_1 gpc1_1_490(
      {stage24[13]},
      {stage24[86]}
   );
   gpc1_1 gpc1_1_491(
      {stage24[14]},
      {stage24[87]}
   );
   gpc1_1 gpc1_1_492(
      {stage24[15]},
      {stage24[88]}
   );
   gpc606_5 gpc606_5_493(
      {stage24[16], stage24[17], stage24[18], stage24[19], stage24[20], stage24[21]},
      {stage26[0], stage26[1], stage26[2], stage26[3], stage26[4], stage26[5]},
      {stage28[64], stage27[67], stage26[68], stage25[74], stage24[89]}
   );
   gpc615_5 gpc615_5_494(
      {stage24[22], stage24[23], stage24[24], stage24[25], stage24[26]},
      {stage25[18]},
      {stage26[6], stage26[7], stage26[8], stage26[9], stage26[10], stage26[11]},
      {stage28[65], stage27[68], stage26[69], stage25[75], stage24[90]}
   );
   gpc615_5 gpc615_5_495(
      {stage24[27], stage24[28], stage24[29], stage24[30], stage24[31]},
      {stage25[19]},
      {stage26[12], stage26[13], stage26[14], stage26[15], stage26[16], stage26[17]},
      {stage28[66], stage27[69], stage26[70], stage25[76], stage24[91]}
   );
   gpc615_5 gpc615_5_496(
      {stage24[32], stage24[33], stage24[34], stage24[35], stage24[36]},
      {stage25[20]},
      {stage26[18], stage26[19], stage26[20], stage26[21], stage26[22], stage26[23]},
      {stage28[67], stage27[70], stage26[71], stage25[77], stage24[92]}
   );
   gpc615_5 gpc615_5_497(
      {stage24[37], stage24[38], stage24[39], stage24[40], stage24[41]},
      {stage25[21]},
      {stage26[24], stage26[25], stage26[26], stage26[27], stage26[28], stage26[29]},
      {stage28[68], stage27[71], stage26[72], stage25[78], stage24[93]}
   );
   gpc615_5 gpc615_5_498(
      {stage24[42], stage24[43], stage24[44], stage24[45], stage24[46]},
      {stage25[22]},
      {stage26[30], stage26[31], stage26[32], stage26[33], stage26[34], stage26[35]},
      {stage28[69], stage27[72], stage26[73], stage25[79], stage24[94]}
   );
   gpc615_5 gpc615_5_499(
      {stage24[47], stage24[48], stage24[49], stage24[50], stage24[51]},
      {stage25[23]},
      {stage26[36], stage26[37], stage26[38], stage26[39], stage26[40], stage26[41]},
      {stage28[70], stage27[73], stage26[74], stage25[80], stage24[95]}
   );
   gpc135_4 gpc135_4_500(
      {stage24[52], stage24[53], stage24[54], stage24[55], stage24[56]},
      {stage25[24], stage25[25], stage25[26]},
      {stage26[42]},
      {stage27[74], stage26[75], stage25[81], stage24[96]}
   );
   gpc207_4 gpc207_4_501(
      {stage24[57], stage24[58], stage24[59], stage24[60], stage24[61], stage24[62], stage24[63]},
      {stage26[43], stage26[44]},
      {stage27[75], stage26[76], stage25[82], stage24[97]}
   );
   gpc1_1 gpc1_1_502(
      {stage25[27]},
      {stage25[83]}
   );
   gpc1_1 gpc1_1_503(
      {stage25[28]},
      {stage25[84]}
   );
   gpc1_1 gpc1_1_504(
      {stage25[29]},
      {stage25[85]}
   );
   gpc1_1 gpc1_1_505(
      {stage25[30]},
      {stage25[86]}
   );
   gpc1_1 gpc1_1_506(
      {stage25[31]},
      {stage25[87]}
   );
   gpc1_1 gpc1_1_507(
      {stage25[32]},
      {stage25[88]}
   );
   gpc1_1 gpc1_1_508(
      {stage25[33]},
      {stage25[89]}
   );
   gpc1_1 gpc1_1_509(
      {stage25[34]},
      {stage25[90]}
   );
   gpc1_1 gpc1_1_510(
      {stage25[35]},
      {stage25[91]}
   );
   gpc1_1 gpc1_1_511(
      {stage25[36]},
      {stage25[92]}
   );
   gpc606_5 gpc606_5_512(
      {stage25[37], stage25[38], stage25[39], stage25[40], stage25[41], stage25[42]},
      {stage27[0], stage27[1], stage27[2], stage27[3], stage27[4], stage27[5]},
      {stage29[64], stage28[71], stage27[76], stage26[77], stage25[93]}
   );
   gpc606_5 gpc606_5_513(
      {stage25[43], stage25[44], stage25[45], stage25[46], stage25[47], stage25[48]},
      {stage27[6], stage27[7], stage27[8], stage27[9], stage27[10], stage27[11]},
      {stage29[65], stage28[72], stage27[77], stage26[78], stage25[94]}
   );
   gpc606_5 gpc606_5_514(
      {stage25[49], stage25[50], stage25[51], stage25[52], stage25[53], stage25[54]},
      {stage27[12], stage27[13], stage27[14], stage27[15], stage27[16], stage27[17]},
      {stage29[66], stage28[73], stage27[78], stage26[79], stage25[95]}
   );
   gpc606_5 gpc606_5_515(
      {stage25[55], stage25[56], stage25[57], stage25[58], stage25[59], stage25[60]},
      {stage27[18], stage27[19], stage27[20], stage27[21], stage27[22], stage27[23]},
      {stage29[67], stage28[74], stage27[79], stage26[80], stage25[96]}
   );
   gpc1343_5 gpc1343_5_516(
      {stage25[61], stage25[62], stage25[63]},
      {stage26[45], stage26[46], stage26[47], stage26[48]},
      {stage27[24], stage27[25], stage27[26]},
      {stage28[0]},
      {stage29[68], stage28[75], stage27[80], stage26[81], stage25[97]}
   );
   gpc1_1 gpc1_1_517(
      {stage26[49]},
      {stage26[82]}
   );
   gpc1_1 gpc1_1_518(
      {stage26[50]},
      {stage26[83]}
   );
   gpc1_1 gpc1_1_519(
      {stage26[51]},
      {stage26[84]}
   );
   gpc606_5 gpc606_5_520(
      {stage26[52], stage26[53], stage26[54], stage26[55], stage26[56], stage26[57]},
      {stage28[1], stage28[2], stage28[3], stage28[4], stage28[5], stage28[6]},
      {stage30[64], stage29[69], stage28[76], stage27[81], stage26[85]}
   );
   gpc606_5 gpc606_5_521(
      {stage26[58], stage26[59], stage26[60], stage26[61], stage26[62], stage26[63]},
      {stage28[7], stage28[8], stage28[9], stage28[10], stage28[11], stage28[12]},
      {stage30[65], stage29[70], stage28[77], stage27[82], stage26[86]}
   );
   gpc1_1 gpc1_1_522(
      {stage27[27]},
      {stage27[83]}
   );
   gpc1_1 gpc1_1_523(
      {stage27[28]},
      {stage27[84]}
   );
   gpc1_1 gpc1_1_524(
      {stage27[29]},
      {stage27[85]}
   );
   gpc1_1 gpc1_1_525(
      {stage27[30]},
      {stage27[86]}
   );
   gpc1_1 gpc1_1_526(
      {stage27[31]},
      {stage27[87]}
   );
   gpc1_1 gpc1_1_527(
      {stage27[32]},
      {stage27[88]}
   );
   gpc1_1 gpc1_1_528(
      {stage27[33]},
      {stage27[89]}
   );
   gpc1_1 gpc1_1_529(
      {stage27[34]},
      {stage27[90]}
   );
   gpc1_1 gpc1_1_530(
      {stage27[35]},
      {stage27[91]}
   );
   gpc1_1 gpc1_1_531(
      {stage27[36]},
      {stage27[92]}
   );
   gpc1_1 gpc1_1_532(
      {stage27[37]},
      {stage27[93]}
   );
   gpc1_1 gpc1_1_533(
      {stage27[38]},
      {stage27[94]}
   );
   gpc1_1 gpc1_1_534(
      {stage27[39]},
      {stage27[95]}
   );
   gpc1_1 gpc1_1_535(
      {stage27[40]},
      {stage27[96]}
   );
   gpc1_1 gpc1_1_536(
      {stage27[41]},
      {stage27[97]}
   );
   gpc1_1 gpc1_1_537(
      {stage27[42]},
      {stage27[98]}
   );
   gpc1_1 gpc1_1_538(
      {stage27[43]},
      {stage27[99]}
   );
   gpc615_5 gpc615_5_539(
      {stage27[44], stage27[45], stage27[46], stage27[47], stage27[48]},
      {stage28[13]},
      {stage29[0], stage29[1], stage29[2], stage29[3], stage29[4], stage29[5]},
      {stage31[64], stage30[66], stage29[71], stage28[78], stage27[100]}
   );
   gpc615_5 gpc615_5_540(
      {stage27[49], stage27[50], stage27[51], stage27[52], stage27[53]},
      {stage28[14]},
      {stage29[6], stage29[7], stage29[8], stage29[9], stage29[10], stage29[11]},
      {stage31[65], stage30[67], stage29[72], stage28[79], stage27[101]}
   );
   gpc615_5 gpc615_5_541(
      {stage27[54], stage27[55], stage27[56], stage27[57], stage27[58]},
      {stage28[15]},
      {stage29[12], stage29[13], stage29[14], stage29[15], stage29[16], stage29[17]},
      {stage31[66], stage30[68], stage29[73], stage28[80], stage27[102]}
   );
   gpc615_5 gpc615_5_542(
      {stage27[59], stage27[60], stage27[61], stage27[62], stage27[63]},
      {stage28[16]},
      {stage29[18], stage29[19], stage29[20], stage29[21], stage29[22], stage29[23]},
      {stage31[67], stage30[69], stage29[74], stage28[81], stage27[103]}
   );
   gpc606_5 gpc606_5_543(
      {stage28[17], stage28[18], stage28[19], stage28[20], stage28[21], stage28[22]},
      {stage30[0], stage30[1], stage30[2], stage30[3], stage30[4], stage30[5]},
      {stage32[64], stage31[68], stage30[70], stage29[75], stage28[82]}
   );
   gpc606_5 gpc606_5_544(
      {stage28[23], stage28[24], stage28[25], stage28[26], stage28[27], stage28[28]},
      {stage30[6], stage30[7], stage30[8], stage30[9], stage30[10], stage30[11]},
      {stage32[65], stage31[69], stage30[71], stage29[76], stage28[83]}
   );
   gpc606_5 gpc606_5_545(
      {stage28[29], stage28[30], stage28[31], stage28[32], stage28[33], stage28[34]},
      {stage30[12], stage30[13], stage30[14], stage30[15], stage30[16], stage30[17]},
      {stage32[66], stage31[70], stage30[72], stage29[77], stage28[84]}
   );
   gpc606_5 gpc606_5_546(
      {stage28[35], stage28[36], stage28[37], stage28[38], stage28[39], stage28[40]},
      {stage30[18], stage30[19], stage30[20], stage30[21], stage30[22], stage30[23]},
      {stage32[67], stage31[71], stage30[73], stage29[78], stage28[85]}
   );
   gpc606_5 gpc606_5_547(
      {stage28[41], stage28[42], stage28[43], stage28[44], stage28[45], stage28[46]},
      {stage30[24], stage30[25], stage30[26], stage30[27], stage30[28], stage30[29]},
      {stage32[68], stage31[72], stage30[74], stage29[79], stage28[86]}
   );
   gpc606_5 gpc606_5_548(
      {stage28[47], stage28[48], stage28[49], stage28[50], stage28[51], stage28[52]},
      {stage30[30], stage30[31], stage30[32], stage30[33], stage30[34], stage30[35]},
      {stage32[69], stage31[73], stage30[75], stage29[80], stage28[87]}
   );
   gpc606_5 gpc606_5_549(
      {stage28[53], stage28[54], stage28[55], stage28[56], stage28[57], stage28[58]},
      {stage30[36], stage30[37], stage30[38], stage30[39], stage30[40], stage30[41]},
      {stage32[70], stage31[74], stage30[76], stage29[81], stage28[88]}
   );
   gpc606_5 gpc606_5_550(
      {stage28[59], stage28[60], stage28[61], stage28[62], stage28[63], 1'h0},
      {stage30[42], stage30[43], stage30[44], stage30[45], stage30[46], stage30[47]},
      {stage32[71], stage31[75], stage30[77], stage29[82], stage28[89]}
   );
   gpc1_1 gpc1_1_551(
      {stage29[24]},
      {stage29[83]}
   );
   gpc1_1 gpc1_1_552(
      {stage29[25]},
      {stage29[84]}
   );
   gpc1_1 gpc1_1_553(
      {stage29[26]},
      {stage29[85]}
   );
   gpc1_1 gpc1_1_554(
      {stage29[27]},
      {stage29[86]}
   );
   gpc1_1 gpc1_1_555(
      {stage29[28]},
      {stage29[87]}
   );
   gpc606_5 gpc606_5_556(
      {stage29[29], stage29[30], stage29[31], stage29[32], stage29[33], stage29[34]},
      {stage31[0], stage31[1], stage31[2], stage31[3], stage31[4], stage31[5]},
      {stage33[64], stage32[72], stage31[76], stage30[78], stage29[88]}
   );
   gpc606_5 gpc606_5_557(
      {stage29[35], stage29[36], stage29[37], stage29[38], stage29[39], stage29[40]},
      {stage31[6], stage31[7], stage31[8], stage31[9], stage31[10], stage31[11]},
      {stage33[65], stage32[73], stage31[77], stage30[79], stage29[89]}
   );
   gpc606_5 gpc606_5_558(
      {stage29[41], stage29[42], stage29[43], stage29[44], stage29[45], stage29[46]},
      {stage31[12], stage31[13], stage31[14], stage31[15], stage31[16], stage31[17]},
      {stage33[66], stage32[74], stage31[78], stage30[80], stage29[90]}
   );
   gpc606_5 gpc606_5_559(
      {stage29[47], stage29[48], stage29[49], stage29[50], stage29[51], stage29[52]},
      {stage31[18], stage31[19], stage31[20], stage31[21], stage31[22], stage31[23]},
      {stage33[67], stage32[75], stage31[79], stage30[81], stage29[91]}
   );
   gpc606_5 gpc606_5_560(
      {stage29[53], stage29[54], stage29[55], stage29[56], stage29[57], stage29[58]},
      {stage31[24], stage31[25], stage31[26], stage31[27], stage31[28], stage31[29]},
      {stage33[68], stage32[76], stage31[80], stage30[82], stage29[92]}
   );
   gpc615_5 gpc615_5_561(
      {stage29[59], stage29[60], stage29[61], stage29[62], stage29[63]},
      {stage30[48]},
      {stage31[30], stage31[31], stage31[32], stage31[33], stage31[34], stage31[35]},
      {stage33[69], stage32[77], stage31[81], stage30[83], stage29[93]}
   );
   gpc1_1 gpc1_1_562(
      {stage30[49]},
      {stage30[84]}
   );
   gpc1_1 gpc1_1_563(
      {stage30[50]},
      {stage30[85]}
   );
   gpc1_1 gpc1_1_564(
      {stage30[51]},
      {stage30[86]}
   );
   gpc1_1 gpc1_1_565(
      {stage30[52]},
      {stage30[87]}
   );
   gpc1_1 gpc1_1_566(
      {stage30[53]},
      {stage30[88]}
   );
   gpc1_1 gpc1_1_567(
      {stage30[54]},
      {stage30[89]}
   );
   gpc1_1 gpc1_1_568(
      {stage30[55]},
      {stage30[90]}
   );
   gpc1_1 gpc1_1_569(
      {stage30[56]},
      {stage30[91]}
   );
   gpc1_1 gpc1_1_570(
      {stage30[57]},
      {stage30[92]}
   );
   gpc606_5 gpc606_5_571(
      {stage30[58], stage30[59], stage30[60], stage30[61], stage30[62], stage30[63]},
      {stage32[0], stage32[1], stage32[2], stage32[3], stage32[4], stage32[5]},
      {stage34[64], stage33[70], stage32[78], stage31[82], stage30[93]}
   );
   gpc1_1 gpc1_1_572(
      {stage31[36]},
      {stage31[83]}
   );
   gpc1_1 gpc1_1_573(
      {stage31[37]},
      {stage31[84]}
   );
   gpc1_1 gpc1_1_574(
      {stage31[38]},
      {stage31[85]}
   );
   gpc615_5 gpc615_5_575(
      {stage31[39], stage31[40], stage31[41], stage31[42], stage31[43]},
      {stage32[6]},
      {stage33[0], stage33[1], stage33[2], stage33[3], stage33[4], stage33[5]},
      {stage35[64], stage34[65], stage33[71], stage32[79], stage31[86]}
   );
   gpc615_5 gpc615_5_576(
      {stage31[44], stage31[45], stage31[46], stage31[47], stage31[48]},
      {stage32[7]},
      {stage33[6], stage33[7], stage33[8], stage33[9], stage33[10], stage33[11]},
      {stage35[65], stage34[66], stage33[72], stage32[80], stage31[87]}
   );
   gpc615_5 gpc615_5_577(
      {stage31[49], stage31[50], stage31[51], stage31[52], stage31[53]},
      {stage32[8]},
      {stage33[12], stage33[13], stage33[14], stage33[15], stage33[16], stage33[17]},
      {stage35[66], stage34[67], stage33[73], stage32[81], stage31[88]}
   );
   gpc615_5 gpc615_5_578(
      {stage31[54], stage31[55], stage31[56], stage31[57], stage31[58]},
      {stage32[9]},
      {stage33[18], stage33[19], stage33[20], stage33[21], stage33[22], stage33[23]},
      {stage35[67], stage34[68], stage33[74], stage32[82], stage31[89]}
   );
   gpc615_5 gpc615_5_579(
      {stage31[59], stage31[60], stage31[61], stage31[62], stage31[63]},
      {stage32[10]},
      {stage33[24], stage33[25], stage33[26], stage33[27], stage33[28], stage33[29]},
      {stage35[68], stage34[69], stage33[75], stage32[83], stage31[90]}
   );
   gpc1_1 gpc1_1_580(
      {stage32[11]},
      {stage32[84]}
   );
   gpc1_1 gpc1_1_581(
      {stage32[12]},
      {stage32[85]}
   );
   gpc1_1 gpc1_1_582(
      {stage32[13]},
      {stage32[86]}
   );
   gpc1_1 gpc1_1_583(
      {stage32[14]},
      {stage32[87]}
   );
   gpc1_1 gpc1_1_584(
      {stage32[15]},
      {stage32[88]}
   );
   gpc606_5 gpc606_5_585(
      {stage32[16], stage32[17], stage32[18], stage32[19], stage32[20], stage32[21]},
      {stage34[0], stage34[1], stage34[2], stage34[3], stage34[4], stage34[5]},
      {stage36[64], stage35[69], stage34[70], stage33[76], stage32[89]}
   );
   gpc606_5 gpc606_5_586(
      {stage32[22], stage32[23], stage32[24], stage32[25], stage32[26], stage32[27]},
      {stage34[6], stage34[7], stage34[8], stage34[9], stage34[10], stage34[11]},
      {stage36[65], stage35[70], stage34[71], stage33[77], stage32[90]}
   );
   gpc606_5 gpc606_5_587(
      {stage32[28], stage32[29], stage32[30], stage32[31], stage32[32], stage32[33]},
      {stage34[12], stage34[13], stage34[14], stage34[15], stage34[16], stage34[17]},
      {stage36[66], stage35[71], stage34[72], stage33[78], stage32[91]}
   );
   gpc606_5 gpc606_5_588(
      {stage32[34], stage32[35], stage32[36], stage32[37], stage32[38], stage32[39]},
      {stage34[18], stage34[19], stage34[20], stage34[21], stage34[22], stage34[23]},
      {stage36[67], stage35[72], stage34[73], stage33[79], stage32[92]}
   );
   gpc606_5 gpc606_5_589(
      {stage32[40], stage32[41], stage32[42], stage32[43], stage32[44], stage32[45]},
      {stage34[24], stage34[25], stage34[26], stage34[27], stage34[28], stage34[29]},
      {stage36[68], stage35[73], stage34[74], stage33[80], stage32[93]}
   );
   gpc606_5 gpc606_5_590(
      {stage32[46], stage32[47], stage32[48], stage32[49], stage32[50], stage32[51]},
      {stage34[30], stage34[31], stage34[32], stage34[33], stage34[34], stage34[35]},
      {stage36[69], stage35[74], stage34[75], stage33[81], stage32[94]}
   );
   gpc606_5 gpc606_5_591(
      {stage32[52], stage32[53], stage32[54], stage32[55], stage32[56], stage32[57]},
      {stage34[36], stage34[37], stage34[38], stage34[39], stage34[40], stage34[41]},
      {stage36[70], stage35[75], stage34[76], stage33[82], stage32[95]}
   );
   gpc606_5 gpc606_5_592(
      {stage32[58], stage32[59], stage32[60], stage32[61], stage32[62], stage32[63]},
      {stage34[42], stage34[43], stage34[44], stage34[45], stage34[46], stage34[47]},
      {stage36[71], stage35[76], stage34[77], stage33[83], stage32[96]}
   );
   gpc606_5 gpc606_5_593(
      {stage33[30], stage33[31], stage33[32], stage33[33], stage33[34], stage33[35]},
      {stage35[0], stage35[1], stage35[2], stage35[3], stage35[4], stage35[5]},
      {stage37[64], stage36[72], stage35[77], stage34[78], stage33[84]}
   );
   gpc606_5 gpc606_5_594(
      {stage33[36], stage33[37], stage33[38], stage33[39], stage33[40], stage33[41]},
      {stage35[6], stage35[7], stage35[8], stage35[9], stage35[10], stage35[11]},
      {stage37[65], stage36[73], stage35[78], stage34[79], stage33[85]}
   );
   gpc606_5 gpc606_5_595(
      {stage33[42], stage33[43], stage33[44], stage33[45], stage33[46], stage33[47]},
      {stage35[12], stage35[13], stage35[14], stage35[15], stage35[16], stage35[17]},
      {stage37[66], stage36[74], stage35[79], stage34[80], stage33[86]}
   );
   gpc606_5 gpc606_5_596(
      {stage33[48], stage33[49], stage33[50], stage33[51], stage33[52], stage33[53]},
      {stage35[18], stage35[19], stage35[20], stage35[21], stage35[22], stage35[23]},
      {stage37[67], stage36[75], stage35[80], stage34[81], stage33[87]}
   );
   gpc606_5 gpc606_5_597(
      {stage33[54], stage33[55], stage33[56], stage33[57], stage33[58], stage33[59]},
      {stage35[24], stage35[25], stage35[26], stage35[27], stage35[28], stage35[29]},
      {stage37[68], stage36[76], stage35[81], stage34[82], stage33[88]}
   );
   gpc606_5 gpc606_5_598(
      {stage33[60], stage33[61], stage33[62], stage33[63], 1'h0, 1'h0},
      {stage35[30], stage35[31], stage35[32], stage35[33], stage35[34], stage35[35]},
      {stage37[69], stage36[77], stage35[82], stage34[83], stage33[89]}
   );
   gpc1_1 gpc1_1_599(
      {stage34[48]},
      {stage34[84]}
   );
   gpc615_5 gpc615_5_600(
      {stage34[49], stage34[50], stage34[51], stage34[52], stage34[53]},
      {stage35[36]},
      {stage36[0], stage36[1], stage36[2], stage36[3], stage36[4], stage36[5]},
      {stage38[64], stage37[70], stage36[78], stage35[83], stage34[85]}
   );
   gpc615_5 gpc615_5_601(
      {stage34[54], stage34[55], stage34[56], stage34[57], stage34[58]},
      {stage35[37]},
      {stage36[6], stage36[7], stage36[8], stage36[9], stage36[10], stage36[11]},
      {stage38[65], stage37[71], stage36[79], stage35[84], stage34[86]}
   );
   gpc615_5 gpc615_5_602(
      {stage34[59], stage34[60], stage34[61], stage34[62], stage34[63]},
      {stage35[38]},
      {stage36[12], stage36[13], stage36[14], stage36[15], stage36[16], stage36[17]},
      {stage38[66], stage37[72], stage36[80], stage35[85], stage34[87]}
   );
   gpc615_5 gpc615_5_603(
      {stage35[39], stage35[40], stage35[41], stage35[42], stage35[43]},
      {stage36[18]},
      {stage37[0], stage37[1], stage37[2], stage37[3], stage37[4], stage37[5]},
      {stage39[64], stage38[67], stage37[73], stage36[81], stage35[86]}
   );
   gpc615_5 gpc615_5_604(
      {stage35[44], stage35[45], stage35[46], stage35[47], stage35[48]},
      {stage36[19]},
      {stage37[6], stage37[7], stage37[8], stage37[9], stage37[10], stage37[11]},
      {stage39[65], stage38[68], stage37[74], stage36[82], stage35[87]}
   );
   gpc615_5 gpc615_5_605(
      {stage35[49], stage35[50], stage35[51], stage35[52], stage35[53]},
      {stage36[20]},
      {stage37[12], stage37[13], stage37[14], stage37[15], stage37[16], stage37[17]},
      {stage39[66], stage38[69], stage37[75], stage36[83], stage35[88]}
   );
   gpc615_5 gpc615_5_606(
      {stage35[54], stage35[55], stage35[56], stage35[57], stage35[58]},
      {stage36[21]},
      {stage37[18], stage37[19], stage37[20], stage37[21], stage37[22], stage37[23]},
      {stage39[67], stage38[70], stage37[76], stage36[84], stage35[89]}
   );
   gpc615_5 gpc615_5_607(
      {stage35[59], stage35[60], stage35[61], stage35[62], stage35[63]},
      {stage36[22]},
      {stage37[24], stage37[25], stage37[26], stage37[27], stage37[28], stage37[29]},
      {stage39[68], stage38[71], stage37[77], stage36[85], stage35[90]}
   );
   gpc1_1 gpc1_1_608(
      {stage36[23]},
      {stage36[86]}
   );
   gpc1_1 gpc1_1_609(
      {stage36[24]},
      {stage36[87]}
   );
   gpc1_1 gpc1_1_610(
      {stage36[25]},
      {stage36[88]}
   );
   gpc1_1 gpc1_1_611(
      {stage36[26]},
      {stage36[89]}
   );
   gpc1_1 gpc1_1_612(
      {stage36[27]},
      {stage36[90]}
   );
   gpc1_1 gpc1_1_613(
      {stage36[28]},
      {stage36[91]}
   );
   gpc1_1 gpc1_1_614(
      {stage36[29]},
      {stage36[92]}
   );
   gpc1_1 gpc1_1_615(
      {stage36[30]},
      {stage36[93]}
   );
   gpc1_1 gpc1_1_616(
      {stage36[31]},
      {stage36[94]}
   );
   gpc1_1 gpc1_1_617(
      {stage36[32]},
      {stage36[95]}
   );
   gpc1_1 gpc1_1_618(
      {stage36[33]},
      {stage36[96]}
   );
   gpc1_1 gpc1_1_619(
      {stage36[34]},
      {stage36[97]}
   );
   gpc1_1 gpc1_1_620(
      {stage36[35]},
      {stage36[98]}
   );
   gpc1_1 gpc1_1_621(
      {stage36[36]},
      {stage36[99]}
   );
   gpc1_1 gpc1_1_622(
      {stage36[37]},
      {stage36[100]}
   );
   gpc1_1 gpc1_1_623(
      {stage36[38]},
      {stage36[101]}
   );
   gpc1_1 gpc1_1_624(
      {stage36[39]},
      {stage36[102]}
   );
   gpc606_5 gpc606_5_625(
      {stage36[40], stage36[41], stage36[42], stage36[43], stage36[44], stage36[45]},
      {stage38[0], stage38[1], stage38[2], stage38[3], stage38[4], stage38[5]},
      {stage40[64], stage39[69], stage38[72], stage37[78], stage36[103]}
   );
   gpc606_5 gpc606_5_626(
      {stage36[46], stage36[47], stage36[48], stage36[49], stage36[50], stage36[51]},
      {stage38[6], stage38[7], stage38[8], stage38[9], stage38[10], stage38[11]},
      {stage40[65], stage39[70], stage38[73], stage37[79], stage36[104]}
   );
   gpc606_5 gpc606_5_627(
      {stage36[52], stage36[53], stage36[54], stage36[55], stage36[56], stage36[57]},
      {stage38[12], stage38[13], stage38[14], stage38[15], stage38[16], stage38[17]},
      {stage40[66], stage39[71], stage38[74], stage37[80], stage36[105]}
   );
   gpc606_5 gpc606_5_628(
      {stage36[58], stage36[59], stage36[60], stage36[61], stage36[62], stage36[63]},
      {stage38[18], stage38[19], stage38[20], stage38[21], stage38[22], stage38[23]},
      {stage40[67], stage39[72], stage38[75], stage37[81], stage36[106]}
   );
   gpc1_1 gpc1_1_629(
      {stage37[30]},
      {stage37[82]}
   );
   gpc1_1 gpc1_1_630(
      {stage37[31]},
      {stage37[83]}
   );
   gpc1_1 gpc1_1_631(
      {stage37[32]},
      {stage37[84]}
   );
   gpc1_1 gpc1_1_632(
      {stage37[33]},
      {stage37[85]}
   );
   gpc1_1 gpc1_1_633(
      {stage37[34]},
      {stage37[86]}
   );
   gpc1_1 gpc1_1_634(
      {stage37[35]},
      {stage37[87]}
   );
   gpc1_1 gpc1_1_635(
      {stage37[36]},
      {stage37[88]}
   );
   gpc1_1 gpc1_1_636(
      {stage37[37]},
      {stage37[89]}
   );
   gpc1_1 gpc1_1_637(
      {stage37[38]},
      {stage37[90]}
   );
   gpc1_1 gpc1_1_638(
      {stage37[39]},
      {stage37[91]}
   );
   gpc606_5 gpc606_5_639(
      {stage37[40], stage37[41], stage37[42], stage37[43], stage37[44], stage37[45]},
      {stage39[0], stage39[1], stage39[2], stage39[3], stage39[4], stage39[5]},
      {stage41[64], stage40[68], stage39[73], stage38[76], stage37[92]}
   );
   gpc606_5 gpc606_5_640(
      {stage37[46], stage37[47], stage37[48], stage37[49], stage37[50], stage37[51]},
      {stage39[6], stage39[7], stage39[8], stage39[9], stage39[10], stage39[11]},
      {stage41[65], stage40[69], stage39[74], stage38[77], stage37[93]}
   );
   gpc606_5 gpc606_5_641(
      {stage37[52], stage37[53], stage37[54], stage37[55], stage37[56], stage37[57]},
      {stage39[12], stage39[13], stage39[14], stage39[15], stage39[16], stage39[17]},
      {stage41[66], stage40[70], stage39[75], stage38[78], stage37[94]}
   );
   gpc606_5 gpc606_5_642(
      {stage37[58], stage37[59], stage37[60], stage37[61], stage37[62], stage37[63]},
      {stage39[18], stage39[19], stage39[20], stage39[21], stage39[22], stage39[23]},
      {stage41[67], stage40[71], stage39[76], stage38[79], stage37[95]}
   );
   gpc615_5 gpc615_5_643(
      {stage38[24], stage38[25], stage38[26], stage38[27], stage38[28]},
      {stage39[24]},
      {stage40[0], stage40[1], stage40[2], stage40[3], stage40[4], stage40[5]},
      {stage42[64], stage41[68], stage40[72], stage39[77], stage38[80]}
   );
   gpc615_5 gpc615_5_644(
      {stage38[29], stage38[30], stage38[31], stage38[32], stage38[33]},
      {stage39[25]},
      {stage40[6], stage40[7], stage40[8], stage40[9], stage40[10], stage40[11]},
      {stage42[65], stage41[69], stage40[73], stage39[78], stage38[81]}
   );
   gpc615_5 gpc615_5_645(
      {stage38[34], stage38[35], stage38[36], stage38[37], stage38[38]},
      {stage39[26]},
      {stage40[12], stage40[13], stage40[14], stage40[15], stage40[16], stage40[17]},
      {stage42[66], stage41[70], stage40[74], stage39[79], stage38[82]}
   );
   gpc615_5 gpc615_5_646(
      {stage38[39], stage38[40], stage38[41], stage38[42], stage38[43]},
      {stage39[27]},
      {stage40[18], stage40[19], stage40[20], stage40[21], stage40[22], stage40[23]},
      {stage42[67], stage41[71], stage40[75], stage39[80], stage38[83]}
   );
   gpc615_5 gpc615_5_647(
      {stage38[44], stage38[45], stage38[46], stage38[47], stage38[48]},
      {stage39[28]},
      {stage40[24], stage40[25], stage40[26], stage40[27], stage40[28], stage40[29]},
      {stage42[68], stage41[72], stage40[76], stage39[81], stage38[84]}
   );
   gpc615_5 gpc615_5_648(
      {stage38[49], stage38[50], stage38[51], stage38[52], stage38[53]},
      {stage39[29]},
      {stage40[30], stage40[31], stage40[32], stage40[33], stage40[34], stage40[35]},
      {stage42[69], stage41[73], stage40[77], stage39[82], stage38[85]}
   );
   gpc615_5 gpc615_5_649(
      {stage38[54], stage38[55], stage38[56], stage38[57], stage38[58]},
      {stage39[30]},
      {stage40[36], stage40[37], stage40[38], stage40[39], stage40[40], stage40[41]},
      {stage42[70], stage41[74], stage40[78], stage39[83], stage38[86]}
   );
   gpc615_5 gpc615_5_650(
      {stage38[59], stage38[60], stage38[61], stage38[62], stage38[63]},
      {stage39[31]},
      {stage40[42], stage40[43], stage40[44], stage40[45], stage40[46], stage40[47]},
      {stage42[71], stage41[75], stage40[79], stage39[84], stage38[87]}
   );
   gpc1_1 gpc1_1_651(
      {stage39[32]},
      {stage39[85]}
   );
   gpc1_1 gpc1_1_652(
      {stage39[33]},
      {stage39[86]}
   );
   gpc606_5 gpc606_5_653(
      {stage39[34], stage39[35], stage39[36], stage39[37], stage39[38], stage39[39]},
      {stage41[0], stage41[1], stage41[2], stage41[3], stage41[4], stage41[5]},
      {stage43[64], stage42[72], stage41[76], stage40[80], stage39[87]}
   );
   gpc606_5 gpc606_5_654(
      {stage39[40], stage39[41], stage39[42], stage39[43], stage39[44], stage39[45]},
      {stage41[6], stage41[7], stage41[8], stage41[9], stage41[10], stage41[11]},
      {stage43[65], stage42[73], stage41[77], stage40[81], stage39[88]}
   );
   gpc606_5 gpc606_5_655(
      {stage39[46], stage39[47], stage39[48], stage39[49], stage39[50], stage39[51]},
      {stage41[12], stage41[13], stage41[14], stage41[15], stage41[16], stage41[17]},
      {stage43[66], stage42[74], stage41[78], stage40[82], stage39[89]}
   );
   gpc606_5 gpc606_5_656(
      {stage39[52], stage39[53], stage39[54], stage39[55], stage39[56], stage39[57]},
      {stage41[18], stage41[19], stage41[20], stage41[21], stage41[22], stage41[23]},
      {stage43[67], stage42[75], stage41[79], stage40[83], stage39[90]}
   );
   gpc606_5 gpc606_5_657(
      {stage39[58], stage39[59], stage39[60], stage39[61], stage39[62], stage39[63]},
      {stage41[24], stage41[25], stage41[26], stage41[27], stage41[28], stage41[29]},
      {stage43[68], stage42[76], stage41[80], stage40[84], stage39[91]}
   );
   gpc1_1 gpc1_1_658(
      {stage40[48]},
      {stage40[85]}
   );
   gpc1_1 gpc1_1_659(
      {stage40[49]},
      {stage40[86]}
   );
   gpc1_1 gpc1_1_660(
      {stage40[50]},
      {stage40[87]}
   );
   gpc1_1 gpc1_1_661(
      {stage40[51]},
      {stage40[88]}
   );
   gpc1_1 gpc1_1_662(
      {stage40[52]},
      {stage40[89]}
   );
   gpc1_1 gpc1_1_663(
      {stage40[53]},
      {stage40[90]}
   );
   gpc1_1 gpc1_1_664(
      {stage40[54]},
      {stage40[91]}
   );
   gpc1_1 gpc1_1_665(
      {stage40[55]},
      {stage40[92]}
   );
   gpc1_1 gpc1_1_666(
      {stage40[56]},
      {stage40[93]}
   );
   gpc1_1 gpc1_1_667(
      {stage40[57]},
      {stage40[94]}
   );
   gpc1_1 gpc1_1_668(
      {stage40[58]},
      {stage40[95]}
   );
   gpc1_1 gpc1_1_669(
      {stage40[59]},
      {stage40[96]}
   );
   gpc1_1 gpc1_1_670(
      {stage40[60]},
      {stage40[97]}
   );
   gpc1_1 gpc1_1_671(
      {stage40[61]},
      {stage40[98]}
   );
   gpc1_1 gpc1_1_672(
      {stage40[62]},
      {stage40[99]}
   );
   gpc1_1 gpc1_1_673(
      {stage40[63]},
      {stage40[100]}
   );
   gpc1_1 gpc1_1_674(
      {stage41[30]},
      {stage41[81]}
   );
   gpc1_1 gpc1_1_675(
      {stage41[31]},
      {stage41[82]}
   );
   gpc1_1 gpc1_1_676(
      {stage41[32]},
      {stage41[83]}
   );
   gpc1_1 gpc1_1_677(
      {stage41[33]},
      {stage41[84]}
   );
   gpc1_1 gpc1_1_678(
      {stage41[34]},
      {stage41[85]}
   );
   gpc1_1 gpc1_1_679(
      {stage41[35]},
      {stage41[86]}
   );
   gpc1_1 gpc1_1_680(
      {stage41[36]},
      {stage41[87]}
   );
   gpc1_1 gpc1_1_681(
      {stage41[37]},
      {stage41[88]}
   );
   gpc1_1 gpc1_1_682(
      {stage41[38]},
      {stage41[89]}
   );
   gpc1_1 gpc1_1_683(
      {stage41[39]},
      {stage41[90]}
   );
   gpc1_1 gpc1_1_684(
      {stage41[40]},
      {stage41[91]}
   );
   gpc1_1 gpc1_1_685(
      {stage41[41]},
      {stage41[92]}
   );
   gpc1_1 gpc1_1_686(
      {stage41[42]},
      {stage41[93]}
   );
   gpc1_1 gpc1_1_687(
      {stage41[43]},
      {stage41[94]}
   );
   gpc1_1 gpc1_1_688(
      {stage41[44]},
      {stage41[95]}
   );
   gpc1_1 gpc1_1_689(
      {stage41[45]},
      {stage41[96]}
   );
   gpc1_1 gpc1_1_690(
      {stage41[46]},
      {stage41[97]}
   );
   gpc1_1 gpc1_1_691(
      {stage41[47]},
      {stage41[98]}
   );
   gpc1_1 gpc1_1_692(
      {stage41[48]},
      {stage41[99]}
   );
   gpc1_1 gpc1_1_693(
      {stage41[49]},
      {stage41[100]}
   );
   gpc1_1 gpc1_1_694(
      {stage41[50]},
      {stage41[101]}
   );
   gpc1_1 gpc1_1_695(
      {stage41[51]},
      {stage41[102]}
   );
   gpc1_1 gpc1_1_696(
      {stage41[52]},
      {stage41[103]}
   );
   gpc1_1 gpc1_1_697(
      {stage41[53]},
      {stage41[104]}
   );
   gpc1_1 gpc1_1_698(
      {stage41[54]},
      {stage41[105]}
   );
   gpc1_1 gpc1_1_699(
      {stage41[55]},
      {stage41[106]}
   );
   gpc1_1 gpc1_1_700(
      {stage41[56]},
      {stage41[107]}
   );
   gpc1_1 gpc1_1_701(
      {stage41[57]},
      {stage41[108]}
   );
   gpc606_5 gpc606_5_702(
      {stage41[58], stage41[59], stage41[60], stage41[61], stage41[62], stage41[63]},
      {stage43[0], stage43[1], stage43[2], stage43[3], stage43[4], stage43[5]},
      {stage45[64], stage44[64], stage43[69], stage42[77], stage41[109]}
   );
   gpc1_1 gpc1_1_703(
      {stage42[0]},
      {stage42[78]}
   );
   gpc1_1 gpc1_1_704(
      {stage42[1]},
      {stage42[79]}
   );
   gpc1_1 gpc1_1_705(
      {stage42[2]},
      {stage42[80]}
   );
   gpc1_1 gpc1_1_706(
      {stage42[3]},
      {stage42[81]}
   );
   gpc1_1 gpc1_1_707(
      {stage42[4]},
      {stage42[82]}
   );
   gpc1_1 gpc1_1_708(
      {stage42[5]},
      {stage42[83]}
   );
   gpc1_1 gpc1_1_709(
      {stage42[6]},
      {stage42[84]}
   );
   gpc1_1 gpc1_1_710(
      {stage42[7]},
      {stage42[85]}
   );
   gpc1_1 gpc1_1_711(
      {stage42[8]},
      {stage42[86]}
   );
   gpc1_1 gpc1_1_712(
      {stage42[9]},
      {stage42[87]}
   );
   gpc1_1 gpc1_1_713(
      {stage42[10]},
      {stage42[88]}
   );
   gpc1_1 gpc1_1_714(
      {stage42[11]},
      {stage42[89]}
   );
   gpc1_1 gpc1_1_715(
      {stage42[12]},
      {stage42[90]}
   );
   gpc1_1 gpc1_1_716(
      {stage42[13]},
      {stage42[91]}
   );
   gpc1_1 gpc1_1_717(
      {stage42[14]},
      {stage42[92]}
   );
   gpc1_1 gpc1_1_718(
      {stage42[15]},
      {stage42[93]}
   );
   gpc1_1 gpc1_1_719(
      {stage42[16]},
      {stage42[94]}
   );
   gpc1_1 gpc1_1_720(
      {stage42[17]},
      {stage42[95]}
   );
   gpc1_1 gpc1_1_721(
      {stage42[18]},
      {stage42[96]}
   );
   gpc1325_5 gpc1325_5_722(
      {stage42[19], stage42[20], stage42[21], stage42[22], stage42[23]},
      {stage43[6], stage43[7]},
      {stage44[0], stage44[1], stage44[2]},
      {stage45[0]},
      {stage46[64], stage45[65], stage44[65], stage43[70], stage42[97]}
   );
   gpc1325_5 gpc1325_5_723(
      {stage42[24], stage42[25], stage42[26], stage42[27], stage42[28]},
      {stage43[8], stage43[9]},
      {stage44[3], stage44[4], stage44[5]},
      {stage45[1]},
      {stage46[65], stage45[66], stage44[66], stage43[71], stage42[98]}
   );
   gpc1325_5 gpc1325_5_724(
      {stage42[29], stage42[30], stage42[31], stage42[32], stage42[33]},
      {stage43[10], stage43[11]},
      {stage44[6], stage44[7], stage44[8]},
      {stage45[2]},
      {stage46[66], stage45[67], stage44[67], stage43[72], stage42[99]}
   );
   gpc1325_5 gpc1325_5_725(
      {stage42[34], stage42[35], stage42[36], stage42[37], stage42[38]},
      {stage43[12], stage43[13]},
      {stage44[9], stage44[10], stage44[11]},
      {stage45[3]},
      {stage46[67], stage45[68], stage44[68], stage43[73], stage42[100]}
   );
   gpc1325_5 gpc1325_5_726(
      {stage42[39], stage42[40], stage42[41], stage42[42], stage42[43]},
      {stage43[14], stage43[15]},
      {stage44[12], stage44[13], stage44[14]},
      {stage45[4]},
      {stage46[68], stage45[69], stage44[69], stage43[74], stage42[101]}
   );
   gpc1325_5 gpc1325_5_727(
      {stage42[44], stage42[45], stage42[46], stage42[47], stage42[48]},
      {stage43[16], stage43[17]},
      {stage44[15], stage44[16], stage44[17]},
      {stage45[5]},
      {stage46[69], stage45[70], stage44[70], stage43[75], stage42[102]}
   );
   gpc1325_5 gpc1325_5_728(
      {stage42[49], stage42[50], stage42[51], stage42[52], stage42[53]},
      {stage43[18], stage43[19]},
      {stage44[18], stage44[19], stage44[20]},
      {stage45[6]},
      {stage46[70], stage45[71], stage44[71], stage43[76], stage42[103]}
   );
   gpc1325_5 gpc1325_5_729(
      {stage42[54], stage42[55], stage42[56], stage42[57], stage42[58]},
      {stage43[20], stage43[21]},
      {stage44[21], stage44[22], stage44[23]},
      {stage45[7]},
      {stage46[71], stage45[72], stage44[72], stage43[77], stage42[104]}
   );
   gpc1325_5 gpc1325_5_730(
      {stage42[59], stage42[60], stage42[61], stage42[62], stage42[63]},
      {stage43[22], stage43[23]},
      {stage44[24], stage44[25], stage44[26]},
      {stage45[8]},
      {stage46[72], stage45[73], stage44[73], stage43[78], stage42[105]}
   );
   gpc1_1 gpc1_1_731(
      {stage43[24]},
      {stage43[79]}
   );
   gpc1_1 gpc1_1_732(
      {stage43[25]},
      {stage43[80]}
   );
   gpc1_1 gpc1_1_733(
      {stage43[26]},
      {stage43[81]}
   );
   gpc1_1 gpc1_1_734(
      {stage43[27]},
      {stage43[82]}
   );
   gpc1_1 gpc1_1_735(
      {stage43[28]},
      {stage43[83]}
   );
   gpc1_1 gpc1_1_736(
      {stage43[29]},
      {stage43[84]}
   );
   gpc1_1 gpc1_1_737(
      {stage43[30]},
      {stage43[85]}
   );
   gpc1_1 gpc1_1_738(
      {stage43[31]},
      {stage43[86]}
   );
   gpc1_1 gpc1_1_739(
      {stage43[32]},
      {stage43[87]}
   );
   gpc1_1 gpc1_1_740(
      {stage43[33]},
      {stage43[88]}
   );
   gpc1_1 gpc1_1_741(
      {stage43[34]},
      {stage43[89]}
   );
   gpc1_1 gpc1_1_742(
      {stage43[35]},
      {stage43[90]}
   );
   gpc1_1 gpc1_1_743(
      {stage43[36]},
      {stage43[91]}
   );
   gpc1_1 gpc1_1_744(
      {stage43[37]},
      {stage43[92]}
   );
   gpc1_1 gpc1_1_745(
      {stage43[38]},
      {stage43[93]}
   );
   gpc1_1 gpc1_1_746(
      {stage43[39]},
      {stage43[94]}
   );
   gpc606_5 gpc606_5_747(
      {stage43[40], stage43[41], stage43[42], stage43[43], stage43[44], stage43[45]},
      {stage45[9], stage45[10], stage45[11], stage45[12], stage45[13], stage45[14]},
      {stage47[64], stage46[73], stage45[74], stage44[74], stage43[95]}
   );
   gpc606_5 gpc606_5_748(
      {stage43[46], stage43[47], stage43[48], stage43[49], stage43[50], stage43[51]},
      {stage45[15], stage45[16], stage45[17], stage45[18], stage45[19], stage45[20]},
      {stage47[65], stage46[74], stage45[75], stage44[75], stage43[96]}
   );
   gpc606_5 gpc606_5_749(
      {stage43[52], stage43[53], stage43[54], stage43[55], stage43[56], stage43[57]},
      {stage45[21], stage45[22], stage45[23], stage45[24], stage45[25], stage45[26]},
      {stage47[66], stage46[75], stage45[76], stage44[76], stage43[97]}
   );
   gpc606_5 gpc606_5_750(
      {stage43[58], stage43[59], stage43[60], stage43[61], stage43[62], stage43[63]},
      {stage45[27], stage45[28], stage45[29], stage45[30], stage45[31], stage45[32]},
      {stage47[67], stage46[76], stage45[77], stage44[77], stage43[98]}
   );
   gpc1_1 gpc1_1_751(
      {stage44[27]},
      {stage44[78]}
   );
   gpc606_5 gpc606_5_752(
      {stage44[28], stage44[29], stage44[30], stage44[31], stage44[32], stage44[33]},
      {stage46[0], stage46[1], stage46[2], stage46[3], stage46[4], stage46[5]},
      {stage48[64], stage47[68], stage46[77], stage45[78], stage44[79]}
   );
   gpc606_5 gpc606_5_753(
      {stage44[34], stage44[35], stage44[36], stage44[37], stage44[38], stage44[39]},
      {stage46[6], stage46[7], stage46[8], stage46[9], stage46[10], stage46[11]},
      {stage48[65], stage47[69], stage46[78], stage45[79], stage44[80]}
   );
   gpc606_5 gpc606_5_754(
      {stage44[40], stage44[41], stage44[42], stage44[43], stage44[44], stage44[45]},
      {stage46[12], stage46[13], stage46[14], stage46[15], stage46[16], stage46[17]},
      {stage48[66], stage47[70], stage46[79], stage45[80], stage44[81]}
   );
   gpc606_5 gpc606_5_755(
      {stage44[46], stage44[47], stage44[48], stage44[49], stage44[50], stage44[51]},
      {stage46[18], stage46[19], stage46[20], stage46[21], stage46[22], stage46[23]},
      {stage48[67], stage47[71], stage46[80], stage45[81], stage44[82]}
   );
   gpc606_5 gpc606_5_756(
      {stage44[52], stage44[53], stage44[54], stage44[55], stage44[56], stage44[57]},
      {stage46[24], stage46[25], stage46[26], stage46[27], stage46[28], stage46[29]},
      {stage48[68], stage47[72], stage46[81], stage45[82], stage44[83]}
   );
   gpc606_5 gpc606_5_757(
      {stage44[58], stage44[59], stage44[60], stage44[61], stage44[62], stage44[63]},
      {stage46[30], stage46[31], stage46[32], stage46[33], stage46[34], stage46[35]},
      {stage48[69], stage47[73], stage46[82], stage45[83], stage44[84]}
   );
   gpc1_1 gpc1_1_758(
      {stage45[33]},
      {stage45[84]}
   );
   gpc1_1 gpc1_1_759(
      {stage45[34]},
      {stage45[85]}
   );
   gpc1_1 gpc1_1_760(
      {stage45[35]},
      {stage45[86]}
   );
   gpc623_5 gpc623_5_761(
      {stage45[36], stage45[37], stage45[38]},
      {stage46[36], stage46[37]},
      {stage47[0], stage47[1], stage47[2], stage47[3], stage47[4], stage47[5]},
      {stage49[64], stage48[70], stage47[74], stage46[83], stage45[87]}
   );
   gpc615_5 gpc615_5_762(
      {stage45[39], stage45[40], stage45[41], stage45[42], stage45[43]},
      {stage46[38]},
      {stage47[6], stage47[7], stage47[8], stage47[9], stage47[10], stage47[11]},
      {stage49[65], stage48[71], stage47[75], stage46[84], stage45[88]}
   );
   gpc615_5 gpc615_5_763(
      {stage45[44], stage45[45], stage45[46], stage45[47], stage45[48]},
      {stage46[39]},
      {stage47[12], stage47[13], stage47[14], stage47[15], stage47[16], stage47[17]},
      {stage49[66], stage48[72], stage47[76], stage46[85], stage45[89]}
   );
   gpc615_5 gpc615_5_764(
      {stage45[49], stage45[50], stage45[51], stage45[52], stage45[53]},
      {stage46[40]},
      {stage47[18], stage47[19], stage47[20], stage47[21], stage47[22], stage47[23]},
      {stage49[67], stage48[73], stage47[77], stage46[86], stage45[90]}
   );
   gpc615_5 gpc615_5_765(
      {stage45[54], stage45[55], stage45[56], stage45[57], stage45[58]},
      {stage46[41]},
      {stage47[24], stage47[25], stage47[26], stage47[27], stage47[28], stage47[29]},
      {stage49[68], stage48[74], stage47[78], stage46[87], stage45[91]}
   );
   gpc615_5 gpc615_5_766(
      {stage45[59], stage45[60], stage45[61], stage45[62], stage45[63]},
      {stage46[42]},
      {stage47[30], stage47[31], stage47[32], stage47[33], stage47[34], stage47[35]},
      {stage49[69], stage48[75], stage47[79], stage46[88], stage45[92]}
   );
   gpc1_1 gpc1_1_767(
      {stage46[43]},
      {stage46[89]}
   );
   gpc1_1 gpc1_1_768(
      {stage46[44]},
      {stage46[90]}
   );
   gpc1_1 gpc1_1_769(
      {stage46[45]},
      {stage46[91]}
   );
   gpc1_1 gpc1_1_770(
      {stage46[46]},
      {stage46[92]}
   );
   gpc1_1 gpc1_1_771(
      {stage46[47]},
      {stage46[93]}
   );
   gpc1_1 gpc1_1_772(
      {stage46[48]},
      {stage46[94]}
   );
   gpc1_1 gpc1_1_773(
      {stage46[49]},
      {stage46[95]}
   );
   gpc1_1 gpc1_1_774(
      {stage46[50]},
      {stage46[96]}
   );
   gpc1_1 gpc1_1_775(
      {stage46[51]},
      {stage46[97]}
   );
   gpc1_1 gpc1_1_776(
      {stage46[52]},
      {stage46[98]}
   );
   gpc1_1 gpc1_1_777(
      {stage46[53]},
      {stage46[99]}
   );
   gpc1_1 gpc1_1_778(
      {stage46[54]},
      {stage46[100]}
   );
   gpc1_1 gpc1_1_779(
      {stage46[55]},
      {stage46[101]}
   );
   gpc1_1 gpc1_1_780(
      {stage46[56]},
      {stage46[102]}
   );
   gpc1_1 gpc1_1_781(
      {stage46[57]},
      {stage46[103]}
   );
   gpc1_1 gpc1_1_782(
      {stage46[58]},
      {stage46[104]}
   );
   gpc615_5 gpc615_5_783(
      {stage46[59], stage46[60], stage46[61], stage46[62], stage46[63]},
      {stage47[36]},
      {stage48[0], stage48[1], stage48[2], stage48[3], stage48[4], stage48[5]},
      {stage50[64], stage49[70], stage48[76], stage47[80], stage46[105]}
   );
   gpc1_1 gpc1_1_784(
      {stage47[37]},
      {stage47[81]}
   );
   gpc1_1 gpc1_1_785(
      {stage47[38]},
      {stage47[82]}
   );
   gpc1_1 gpc1_1_786(
      {stage47[39]},
      {stage47[83]}
   );
   gpc1_1 gpc1_1_787(
      {stage47[40]},
      {stage47[84]}
   );
   gpc1_1 gpc1_1_788(
      {stage47[41]},
      {stage47[85]}
   );
   gpc1_1 gpc1_1_789(
      {stage47[42]},
      {stage47[86]}
   );
   gpc615_5 gpc615_5_790(
      {stage47[43], stage47[44], stage47[45], stage47[46], stage47[47]},
      {stage48[6]},
      {stage49[0], stage49[1], stage49[2], stage49[3], stage49[4], stage49[5]},
      {stage51[64], stage50[65], stage49[71], stage48[77], stage47[87]}
   );
   gpc615_5 gpc615_5_791(
      {stage47[48], stage47[49], stage47[50], stage47[51], stage47[52]},
      {stage48[7]},
      {stage49[6], stage49[7], stage49[8], stage49[9], stage49[10], stage49[11]},
      {stage51[65], stage50[66], stage49[72], stage48[78], stage47[88]}
   );
   gpc615_5 gpc615_5_792(
      {stage47[53], stage47[54], stage47[55], stage47[56], stage47[57]},
      {stage48[8]},
      {stage49[12], stage49[13], stage49[14], stage49[15], stage49[16], stage49[17]},
      {stage51[66], stage50[67], stage49[73], stage48[79], stage47[89]}
   );
   gpc1406_5 gpc1406_5_793(
      {stage47[58], stage47[59], stage47[60], stage47[61], stage47[62], stage47[63]},
      {stage49[18], stage49[19], stage49[20], stage49[21]},
      {stage50[0]},
      {stage51[67], stage50[68], stage49[74], stage48[80], stage47[90]}
   );
   gpc1_1 gpc1_1_794(
      {stage48[9]},
      {stage48[81]}
   );
   gpc1_1 gpc1_1_795(
      {stage48[10]},
      {stage48[82]}
   );
   gpc1_1 gpc1_1_796(
      {stage48[11]},
      {stage48[83]}
   );
   gpc1_1 gpc1_1_797(
      {stage48[12]},
      {stage48[84]}
   );
   gpc1_1 gpc1_1_798(
      {stage48[13]},
      {stage48[85]}
   );
   gpc1_1 gpc1_1_799(
      {stage48[14]},
      {stage48[86]}
   );
   gpc1_1 gpc1_1_800(
      {stage48[15]},
      {stage48[87]}
   );
   gpc1_1 gpc1_1_801(
      {stage48[16]},
      {stage48[88]}
   );
   gpc1_1 gpc1_1_802(
      {stage48[17]},
      {stage48[89]}
   );
   gpc1_1 gpc1_1_803(
      {stage48[18]},
      {stage48[90]}
   );
   gpc1_1 gpc1_1_804(
      {stage48[19]},
      {stage48[91]}
   );
   gpc1_1 gpc1_1_805(
      {stage48[20]},
      {stage48[92]}
   );
   gpc1_1 gpc1_1_806(
      {stage48[21]},
      {stage48[93]}
   );
   gpc606_5 gpc606_5_807(
      {stage48[22], stage48[23], stage48[24], stage48[25], stage48[26], stage48[27]},
      {stage50[1], stage50[2], stage50[3], stage50[4], stage50[5], stage50[6]},
      {stage52[64], stage51[68], stage50[69], stage49[75], stage48[94]}
   );
   gpc606_5 gpc606_5_808(
      {stage48[28], stage48[29], stage48[30], stage48[31], stage48[32], stage48[33]},
      {stage50[7], stage50[8], stage50[9], stage50[10], stage50[11], stage50[12]},
      {stage52[65], stage51[69], stage50[70], stage49[76], stage48[95]}
   );
   gpc606_5 gpc606_5_809(
      {stage48[34], stage48[35], stage48[36], stage48[37], stage48[38], stage48[39]},
      {stage50[13], stage50[14], stage50[15], stage50[16], stage50[17], stage50[18]},
      {stage52[66], stage51[70], stage50[71], stage49[77], stage48[96]}
   );
   gpc606_5 gpc606_5_810(
      {stage48[40], stage48[41], stage48[42], stage48[43], stage48[44], stage48[45]},
      {stage50[19], stage50[20], stage50[21], stage50[22], stage50[23], stage50[24]},
      {stage52[67], stage51[71], stage50[72], stage49[78], stage48[97]}
   );
   gpc606_5 gpc606_5_811(
      {stage48[46], stage48[47], stage48[48], stage48[49], stage48[50], stage48[51]},
      {stage50[25], stage50[26], stage50[27], stage50[28], stage50[29], stage50[30]},
      {stage52[68], stage51[72], stage50[73], stage49[79], stage48[98]}
   );
   gpc606_5 gpc606_5_812(
      {stage48[52], stage48[53], stage48[54], stage48[55], stage48[56], stage48[57]},
      {stage50[31], stage50[32], stage50[33], stage50[34], stage50[35], stage50[36]},
      {stage52[69], stage51[73], stage50[74], stage49[80], stage48[99]}
   );
   gpc606_5 gpc606_5_813(
      {stage48[58], stage48[59], stage48[60], stage48[61], stage48[62], stage48[63]},
      {stage50[37], stage50[38], stage50[39], stage50[40], stage50[41], stage50[42]},
      {stage52[70], stage51[74], stage50[75], stage49[81], stage48[100]}
   );
   gpc606_5 gpc606_5_814(
      {stage49[22], stage49[23], stage49[24], stage49[25], stage49[26], stage49[27]},
      {stage51[0], stage51[1], stage51[2], stage51[3], stage51[4], stage51[5]},
      {stage53[64], stage52[71], stage51[75], stage50[76], stage49[82]}
   );
   gpc606_5 gpc606_5_815(
      {stage49[28], stage49[29], stage49[30], stage49[31], stage49[32], stage49[33]},
      {stage51[6], stage51[7], stage51[8], stage51[9], stage51[10], stage51[11]},
      {stage53[65], stage52[72], stage51[76], stage50[77], stage49[83]}
   );
   gpc606_5 gpc606_5_816(
      {stage49[34], stage49[35], stage49[36], stage49[37], stage49[38], stage49[39]},
      {stage51[12], stage51[13], stage51[14], stage51[15], stage51[16], stage51[17]},
      {stage53[66], stage52[73], stage51[77], stage50[78], stage49[84]}
   );
   gpc606_5 gpc606_5_817(
      {stage49[40], stage49[41], stage49[42], stage49[43], stage49[44], stage49[45]},
      {stage51[18], stage51[19], stage51[20], stage51[21], stage51[22], stage51[23]},
      {stage53[67], stage52[74], stage51[78], stage50[79], stage49[85]}
   );
   gpc606_5 gpc606_5_818(
      {stage49[46], stage49[47], stage49[48], stage49[49], stage49[50], stage49[51]},
      {stage51[24], stage51[25], stage51[26], stage51[27], stage51[28], stage51[29]},
      {stage53[68], stage52[75], stage51[79], stage50[80], stage49[86]}
   );
   gpc606_5 gpc606_5_819(
      {stage49[52], stage49[53], stage49[54], stage49[55], stage49[56], stage49[57]},
      {stage51[30], stage51[31], stage51[32], stage51[33], stage51[34], stage51[35]},
      {stage53[69], stage52[76], stage51[80], stage50[81], stage49[87]}
   );
   gpc606_5 gpc606_5_820(
      {stage49[58], stage49[59], stage49[60], stage49[61], stage49[62], stage49[63]},
      {stage51[36], stage51[37], stage51[38], stage51[39], stage51[40], stage51[41]},
      {stage53[70], stage52[77], stage51[81], stage50[82], stage49[88]}
   );
   gpc1_1 gpc1_1_821(
      {stage50[43]},
      {stage50[83]}
   );
   gpc1_1 gpc1_1_822(
      {stage50[44]},
      {stage50[84]}
   );
   gpc1_1 gpc1_1_823(
      {stage50[45]},
      {stage50[85]}
   );
   gpc1_1 gpc1_1_824(
      {stage50[46]},
      {stage50[86]}
   );
   gpc1_1 gpc1_1_825(
      {stage50[47]},
      {stage50[87]}
   );
   gpc1_1 gpc1_1_826(
      {stage50[48]},
      {stage50[88]}
   );
   gpc1_1 gpc1_1_827(
      {stage50[49]},
      {stage50[89]}
   );
   gpc1_1 gpc1_1_828(
      {stage50[50]},
      {stage50[90]}
   );
   gpc1_1 gpc1_1_829(
      {stage50[51]},
      {stage50[91]}
   );
   gpc1_1 gpc1_1_830(
      {stage50[52]},
      {stage50[92]}
   );
   gpc1_1 gpc1_1_831(
      {stage50[53]},
      {stage50[93]}
   );
   gpc615_5 gpc615_5_832(
      {stage50[54], stage50[55], stage50[56], stage50[57], stage50[58]},
      {stage51[42]},
      {stage52[0], stage52[1], stage52[2], stage52[3], stage52[4], stage52[5]},
      {stage54[64], stage53[71], stage52[78], stage51[82], stage50[94]}
   );
   gpc615_5 gpc615_5_833(
      {stage50[59], stage50[60], stage50[61], stage50[62], stage50[63]},
      {stage51[43]},
      {stage52[6], stage52[7], stage52[8], stage52[9], stage52[10], stage52[11]},
      {stage54[65], stage53[72], stage52[79], stage51[83], stage50[95]}
   );
   gpc615_5 gpc615_5_834(
      {stage51[44], stage51[45], stage51[46], stage51[47], stage51[48]},
      {stage52[12]},
      {stage53[0], stage53[1], stage53[2], stage53[3], stage53[4], stage53[5]},
      {stage55[64], stage54[66], stage53[73], stage52[80], stage51[84]}
   );
   gpc615_5 gpc615_5_835(
      {stage51[49], stage51[50], stage51[51], stage51[52], stage51[53]},
      {stage52[13]},
      {stage53[6], stage53[7], stage53[8], stage53[9], stage53[10], stage53[11]},
      {stage55[65], stage54[67], stage53[74], stage52[81], stage51[85]}
   );
   gpc615_5 gpc615_5_836(
      {stage51[54], stage51[55], stage51[56], stage51[57], stage51[58]},
      {stage52[14]},
      {stage53[12], stage53[13], stage53[14], stage53[15], stage53[16], stage53[17]},
      {stage55[66], stage54[68], stage53[75], stage52[82], stage51[86]}
   );
   gpc615_5 gpc615_5_837(
      {stage51[59], stage51[60], stage51[61], stage51[62], stage51[63]},
      {stage52[15]},
      {stage53[18], stage53[19], stage53[20], stage53[21], stage53[22], stage53[23]},
      {stage55[67], stage54[69], stage53[76], stage52[83], stage51[87]}
   );
   gpc606_5 gpc606_5_838(
      {stage52[16], stage52[17], stage52[18], stage52[19], stage52[20], stage52[21]},
      {stage54[0], stage54[1], stage54[2], stage54[3], stage54[4], stage54[5]},
      {stage56[64], stage55[68], stage54[70], stage53[77], stage52[84]}
   );
   gpc606_5 gpc606_5_839(
      {stage52[22], stage52[23], stage52[24], stage52[25], stage52[26], stage52[27]},
      {stage54[6], stage54[7], stage54[8], stage54[9], stage54[10], stage54[11]},
      {stage56[65], stage55[69], stage54[71], stage53[78], stage52[85]}
   );
   gpc606_5 gpc606_5_840(
      {stage52[28], stage52[29], stage52[30], stage52[31], stage52[32], stage52[33]},
      {stage54[12], stage54[13], stage54[14], stage54[15], stage54[16], stage54[17]},
      {stage56[66], stage55[70], stage54[72], stage53[79], stage52[86]}
   );
   gpc606_5 gpc606_5_841(
      {stage52[34], stage52[35], stage52[36], stage52[37], stage52[38], stage52[39]},
      {stage54[18], stage54[19], stage54[20], stage54[21], stage54[22], stage54[23]},
      {stage56[67], stage55[71], stage54[73], stage53[80], stage52[87]}
   );
   gpc606_5 gpc606_5_842(
      {stage52[40], stage52[41], stage52[42], stage52[43], stage52[44], stage52[45]},
      {stage54[24], stage54[25], stage54[26], stage54[27], stage54[28], stage54[29]},
      {stage56[68], stage55[72], stage54[74], stage53[81], stage52[88]}
   );
   gpc606_5 gpc606_5_843(
      {stage52[46], stage52[47], stage52[48], stage52[49], stage52[50], stage52[51]},
      {stage54[30], stage54[31], stage54[32], stage54[33], stage54[34], stage54[35]},
      {stage56[69], stage55[73], stage54[75], stage53[82], stage52[89]}
   );
   gpc606_5 gpc606_5_844(
      {stage52[52], stage52[53], stage52[54], stage52[55], stage52[56], stage52[57]},
      {stage54[36], stage54[37], stage54[38], stage54[39], stage54[40], stage54[41]},
      {stage56[70], stage55[74], stage54[76], stage53[83], stage52[90]}
   );
   gpc606_5 gpc606_5_845(
      {stage52[58], stage52[59], stage52[60], stage52[61], stage52[62], stage52[63]},
      {stage54[42], stage54[43], stage54[44], stage54[45], stage54[46], stage54[47]},
      {stage56[71], stage55[75], stage54[77], stage53[84], stage52[91]}
   );
   gpc1_1 gpc1_1_846(
      {stage53[24]},
      {stage53[85]}
   );
   gpc1_1 gpc1_1_847(
      {stage53[25]},
      {stage53[86]}
   );
   gpc1_1 gpc1_1_848(
      {stage53[26]},
      {stage53[87]}
   );
   gpc1_1 gpc1_1_849(
      {stage53[27]},
      {stage53[88]}
   );
   gpc606_5 gpc606_5_850(
      {stage53[28], stage53[29], stage53[30], stage53[31], stage53[32], stage53[33]},
      {stage55[0], stage55[1], stage55[2], stage55[3], stage55[4], stage55[5]},
      {stage57[64], stage56[72], stage55[76], stage54[78], stage53[89]}
   );
   gpc606_5 gpc606_5_851(
      {stage53[34], stage53[35], stage53[36], stage53[37], stage53[38], stage53[39]},
      {stage55[6], stage55[7], stage55[8], stage55[9], stage55[10], stage55[11]},
      {stage57[65], stage56[73], stage55[77], stage54[79], stage53[90]}
   );
   gpc606_5 gpc606_5_852(
      {stage53[40], stage53[41], stage53[42], stage53[43], stage53[44], stage53[45]},
      {stage55[12], stage55[13], stage55[14], stage55[15], stage55[16], stage55[17]},
      {stage57[66], stage56[74], stage55[78], stage54[80], stage53[91]}
   );
   gpc606_5 gpc606_5_853(
      {stage53[46], stage53[47], stage53[48], stage53[49], stage53[50], stage53[51]},
      {stage55[18], stage55[19], stage55[20], stage55[21], stage55[22], stage55[23]},
      {stage57[67], stage56[75], stage55[79], stage54[81], stage53[92]}
   );
   gpc606_5 gpc606_5_854(
      {stage53[52], stage53[53], stage53[54], stage53[55], stage53[56], stage53[57]},
      {stage55[24], stage55[25], stage55[26], stage55[27], stage55[28], stage55[29]},
      {stage57[68], stage56[76], stage55[80], stage54[82], stage53[93]}
   );
   gpc606_5 gpc606_5_855(
      {stage53[58], stage53[59], stage53[60], stage53[61], stage53[62], stage53[63]},
      {stage55[30], stage55[31], stage55[32], stage55[33], stage55[34], stage55[35]},
      {stage57[69], stage56[77], stage55[81], stage54[83], stage53[94]}
   );
   gpc1_1 gpc1_1_856(
      {stage54[48]},
      {stage54[84]}
   );
   gpc1_1 gpc1_1_857(
      {stage54[49]},
      {stage54[85]}
   );
   gpc1_1 gpc1_1_858(
      {stage54[50]},
      {stage54[86]}
   );
   gpc1_1 gpc1_1_859(
      {stage54[51]},
      {stage54[87]}
   );
   gpc1_1 gpc1_1_860(
      {stage54[52]},
      {stage54[88]}
   );
   gpc1_1 gpc1_1_861(
      {stage54[53]},
      {stage54[89]}
   );
   gpc1_1 gpc1_1_862(
      {stage54[54]},
      {stage54[90]}
   );
   gpc1_1 gpc1_1_863(
      {stage54[55]},
      {stage54[91]}
   );
   gpc1_1 gpc1_1_864(
      {stage54[56]},
      {stage54[92]}
   );
   gpc1_1 gpc1_1_865(
      {stage54[57]},
      {stage54[93]}
   );
   gpc1_1 gpc1_1_866(
      {stage54[58]},
      {stage54[94]}
   );
   gpc1_1 gpc1_1_867(
      {stage54[59]},
      {stage54[95]}
   );
   gpc1_1 gpc1_1_868(
      {stage54[60]},
      {stage54[96]}
   );
   gpc623_5 gpc623_5_869(
      {stage54[61], stage54[62], stage54[63]},
      {stage55[36], stage55[37]},
      {stage56[0], stage56[1], stage56[2], stage56[3], stage56[4], stage56[5]},
      {stage58[64], stage57[70], stage56[78], stage55[82], stage54[97]}
   );
   gpc1_1 gpc1_1_870(
      {stage55[38]},
      {stage55[83]}
   );
   gpc1_1 gpc1_1_871(
      {stage55[39]},
      {stage55[84]}
   );
   gpc1_1 gpc1_1_872(
      {stage55[40]},
      {stage55[85]}
   );
   gpc1_1 gpc1_1_873(
      {stage55[41]},
      {stage55[86]}
   );
   gpc1_1 gpc1_1_874(
      {stage55[42]},
      {stage55[87]}
   );
   gpc1_1 gpc1_1_875(
      {stage55[43]},
      {stage55[88]}
   );
   gpc1_1 gpc1_1_876(
      {stage55[44]},
      {stage55[89]}
   );
   gpc1_1 gpc1_1_877(
      {stage55[45]},
      {stage55[90]}
   );
   gpc606_5 gpc606_5_878(
      {stage55[46], stage55[47], stage55[48], stage55[49], stage55[50], stage55[51]},
      {stage57[0], stage57[1], stage57[2], stage57[3], stage57[4], stage57[5]},
      {stage59[64], stage58[65], stage57[71], stage56[79], stage55[91]}
   );
   gpc606_5 gpc606_5_879(
      {stage55[52], stage55[53], stage55[54], stage55[55], stage55[56], stage55[57]},
      {stage57[6], stage57[7], stage57[8], stage57[9], stage57[10], stage57[11]},
      {stage59[65], stage58[66], stage57[72], stage56[80], stage55[92]}
   );
   gpc606_5 gpc606_5_880(
      {stage55[58], stage55[59], stage55[60], stage55[61], stage55[62], stage55[63]},
      {stage57[12], stage57[13], stage57[14], stage57[15], stage57[16], stage57[17]},
      {stage59[66], stage58[67], stage57[73], stage56[81], stage55[93]}
   );
   gpc1_1 gpc1_1_881(
      {stage56[6]},
      {stage56[82]}
   );
   gpc1_1 gpc1_1_882(
      {stage56[7]},
      {stage56[83]}
   );
   gpc1_1 gpc1_1_883(
      {stage56[8]},
      {stage56[84]}
   );
   gpc1_1 gpc1_1_884(
      {stage56[9]},
      {stage56[85]}
   );
   gpc1_1 gpc1_1_885(
      {stage56[10]},
      {stage56[86]}
   );
   gpc1_1 gpc1_1_886(
      {stage56[11]},
      {stage56[87]}
   );
   gpc1_1 gpc1_1_887(
      {stage56[12]},
      {stage56[88]}
   );
   gpc1_1 gpc1_1_888(
      {stage56[13]},
      {stage56[89]}
   );
   gpc1_1 gpc1_1_889(
      {stage56[14]},
      {stage56[90]}
   );
   gpc1_1 gpc1_1_890(
      {stage56[15]},
      {stage56[91]}
   );
   gpc1_1 gpc1_1_891(
      {stage56[16]},
      {stage56[92]}
   );
   gpc1_1 gpc1_1_892(
      {stage56[17]},
      {stage56[93]}
   );
   gpc1_1 gpc1_1_893(
      {stage56[18]},
      {stage56[94]}
   );
   gpc1_1 gpc1_1_894(
      {stage56[19]},
      {stage56[95]}
   );
   gpc1_1 gpc1_1_895(
      {stage56[20]},
      {stage56[96]}
   );
   gpc1_1 gpc1_1_896(
      {stage56[21]},
      {stage56[97]}
   );
   gpc606_5 gpc606_5_897(
      {stage56[22], stage56[23], stage56[24], stage56[25], stage56[26], stage56[27]},
      {stage58[0], stage58[1], stage58[2], stage58[3], stage58[4], stage58[5]},
      {stage60[64], stage59[67], stage58[68], stage57[74], stage56[98]}
   );
   gpc606_5 gpc606_5_898(
      {stage56[28], stage56[29], stage56[30], stage56[31], stage56[32], stage56[33]},
      {stage58[6], stage58[7], stage58[8], stage58[9], stage58[10], stage58[11]},
      {stage60[65], stage59[68], stage58[69], stage57[75], stage56[99]}
   );
   gpc606_5 gpc606_5_899(
      {stage56[34], stage56[35], stage56[36], stage56[37], stage56[38], stage56[39]},
      {stage58[12], stage58[13], stage58[14], stage58[15], stage58[16], stage58[17]},
      {stage60[66], stage59[69], stage58[70], stage57[76], stage56[100]}
   );
   gpc606_5 gpc606_5_900(
      {stage56[40], stage56[41], stage56[42], stage56[43], stage56[44], stage56[45]},
      {stage58[18], stage58[19], stage58[20], stage58[21], stage58[22], stage58[23]},
      {stage60[67], stage59[70], stage58[71], stage57[77], stage56[101]}
   );
   gpc606_5 gpc606_5_901(
      {stage56[46], stage56[47], stage56[48], stage56[49], stage56[50], stage56[51]},
      {stage58[24], stage58[25], stage58[26], stage58[27], stage58[28], stage58[29]},
      {stage60[68], stage59[71], stage58[72], stage57[78], stage56[102]}
   );
   gpc606_5 gpc606_5_902(
      {stage56[52], stage56[53], stage56[54], stage56[55], stage56[56], stage56[57]},
      {stage58[30], stage58[31], stage58[32], stage58[33], stage58[34], stage58[35]},
      {stage60[69], stage59[72], stage58[73], stage57[79], stage56[103]}
   );
   gpc606_5 gpc606_5_903(
      {stage56[58], stage56[59], stage56[60], stage56[61], stage56[62], stage56[63]},
      {stage58[36], stage58[37], stage58[38], stage58[39], stage58[40], stage58[41]},
      {stage60[70], stage59[73], stage58[74], stage57[80], stage56[104]}
   );
   gpc1_1 gpc1_1_904(
      {stage57[18]},
      {stage57[81]}
   );
   gpc1_1 gpc1_1_905(
      {stage57[19]},
      {stage57[82]}
   );
   gpc1_1 gpc1_1_906(
      {stage57[20]},
      {stage57[83]}
   );
   gpc1_1 gpc1_1_907(
      {stage57[21]},
      {stage57[84]}
   );
   gpc606_5 gpc606_5_908(
      {stage57[22], stage57[23], stage57[24], stage57[25], stage57[26], stage57[27]},
      {stage59[0], stage59[1], stage59[2], stage59[3], stage59[4], stage59[5]},
      {stage61[64], stage60[71], stage59[74], stage58[75], stage57[85]}
   );
   gpc606_5 gpc606_5_909(
      {stage57[28], stage57[29], stage57[30], stage57[31], stage57[32], stage57[33]},
      {stage59[6], stage59[7], stage59[8], stage59[9], stage59[10], stage59[11]},
      {stage61[65], stage60[72], stage59[75], stage58[76], stage57[86]}
   );
   gpc606_5 gpc606_5_910(
      {stage57[34], stage57[35], stage57[36], stage57[37], stage57[38], stage57[39]},
      {stage59[12], stage59[13], stage59[14], stage59[15], stage59[16], stage59[17]},
      {stage61[66], stage60[73], stage59[76], stage58[77], stage57[87]}
   );
   gpc606_5 gpc606_5_911(
      {stage57[40], stage57[41], stage57[42], stage57[43], stage57[44], stage57[45]},
      {stage59[18], stage59[19], stage59[20], stage59[21], stage59[22], stage59[23]},
      {stage61[67], stage60[74], stage59[77], stage58[78], stage57[88]}
   );
   gpc606_5 gpc606_5_912(
      {stage57[46], stage57[47], stage57[48], stage57[49], stage57[50], stage57[51]},
      {stage59[24], stage59[25], stage59[26], stage59[27], stage59[28], stage59[29]},
      {stage61[68], stage60[75], stage59[78], stage58[79], stage57[89]}
   );
   gpc606_5 gpc606_5_913(
      {stage57[52], stage57[53], stage57[54], stage57[55], stage57[56], stage57[57]},
      {stage59[30], stage59[31], stage59[32], stage59[33], stage59[34], stage59[35]},
      {stage61[69], stage60[76], stage59[79], stage58[80], stage57[90]}
   );
   gpc606_5 gpc606_5_914(
      {stage57[58], stage57[59], stage57[60], stage57[61], stage57[62], stage57[63]},
      {stage59[36], stage59[37], stage59[38], stage59[39], stage59[40], stage59[41]},
      {stage61[70], stage60[77], stage59[80], stage58[81], stage57[91]}
   );
   gpc1_1 gpc1_1_915(
      {stage58[42]},
      {stage58[82]}
   );
   gpc1_1 gpc1_1_916(
      {stage58[43]},
      {stage58[83]}
   );
   gpc1_1 gpc1_1_917(
      {stage58[44]},
      {stage58[84]}
   );
   gpc1_1 gpc1_1_918(
      {stage58[45]},
      {stage58[85]}
   );
   gpc1_1 gpc1_1_919(
      {stage58[46]},
      {stage58[86]}
   );
   gpc1_1 gpc1_1_920(
      {stage58[47]},
      {stage58[87]}
   );
   gpc1_1 gpc1_1_921(
      {stage58[48]},
      {stage58[88]}
   );
   gpc1_1 gpc1_1_922(
      {stage58[49]},
      {stage58[89]}
   );
   gpc1_1 gpc1_1_923(
      {stage58[50]},
      {stage58[90]}
   );
   gpc1_1 gpc1_1_924(
      {stage58[51]},
      {stage58[91]}
   );
   gpc1_1 gpc1_1_925(
      {stage58[52]},
      {stage58[92]}
   );
   gpc1_1 gpc1_1_926(
      {stage58[53]},
      {stage58[93]}
   );
   gpc1_1 gpc1_1_927(
      {stage58[54]},
      {stage58[94]}
   );
   gpc1_1 gpc1_1_928(
      {stage58[55]},
      {stage58[95]}
   );
   gpc1_1 gpc1_1_929(
      {stage58[56]},
      {stage58[96]}
   );
   gpc1_1 gpc1_1_930(
      {stage58[57]},
      {stage58[97]}
   );
   gpc606_5 gpc606_5_931(
      {stage58[58], stage58[59], stage58[60], stage58[61], stage58[62], stage58[63]},
      {stage60[0], stage60[1], stage60[2], stage60[3], stage60[4], stage60[5]},
      {stage62[64], stage61[71], stage60[78], stage59[81], stage58[98]}
   );
   gpc1_1 gpc1_1_932(
      {stage59[42]},
      {stage59[82]}
   );
   gpc1_1 gpc1_1_933(
      {stage59[43]},
      {stage59[83]}
   );
   gpc1_1 gpc1_1_934(
      {stage59[44]},
      {stage59[84]}
   );
   gpc1_1 gpc1_1_935(
      {stage59[45]},
      {stage59[85]}
   );
   gpc1_1 gpc1_1_936(
      {stage59[46]},
      {stage59[86]}
   );
   gpc1_1 gpc1_1_937(
      {stage59[47]},
      {stage59[87]}
   );
   gpc1_1 gpc1_1_938(
      {stage59[48]},
      {stage59[88]}
   );
   gpc1_1 gpc1_1_939(
      {stage59[49]},
      {stage59[89]}
   );
   gpc1_1 gpc1_1_940(
      {stage59[50]},
      {stage59[90]}
   );
   gpc1_1 gpc1_1_941(
      {stage59[51]},
      {stage59[91]}
   );
   gpc1_1 gpc1_1_942(
      {stage59[52]},
      {stage59[92]}
   );
   gpc1_1 gpc1_1_943(
      {stage59[53]},
      {stage59[93]}
   );
   gpc1_1 gpc1_1_944(
      {stage59[54]},
      {stage59[94]}
   );
   gpc1_1 gpc1_1_945(
      {stage59[55]},
      {stage59[95]}
   );
   gpc1_1 gpc1_1_946(
      {stage59[56]},
      {stage59[96]}
   );
   gpc1_1 gpc1_1_947(
      {stage59[57]},
      {stage59[97]}
   );
   gpc606_5 gpc606_5_948(
      {stage59[58], stage59[59], stage59[60], stage59[61], stage59[62], stage59[63]},
      {stage61[0], stage61[1], stage61[2], stage61[3], stage61[4], stage61[5]},
      {stage63[64], stage62[65], stage61[72], stage60[79], stage59[98]}
   );
   gpc1_1 gpc1_1_949(
      {stage60[6]},
      {stage60[80]}
   );
   gpc1_1 gpc1_1_950(
      {stage60[7]},
      {stage60[81]}
   );
   gpc1_1 gpc1_1_951(
      {stage60[8]},
      {stage60[82]}
   );
   gpc1_1 gpc1_1_952(
      {stage60[9]},
      {stage60[83]}
   );
   gpc1_1 gpc1_1_953(
      {stage60[10]},
      {stage60[84]}
   );
   gpc1_1 gpc1_1_954(
      {stage60[11]},
      {stage60[85]}
   );
   gpc1_1 gpc1_1_955(
      {stage60[12]},
      {stage60[86]}
   );
   gpc1_1 gpc1_1_956(
      {stage60[13]},
      {stage60[87]}
   );
   gpc1_1 gpc1_1_957(
      {stage60[14]},
      {stage60[88]}
   );
   gpc1_1 gpc1_1_958(
      {stage60[15]},
      {stage60[89]}
   );
   gpc606_5 gpc606_5_959(
      {stage60[16], stage60[17], stage60[18], stage60[19], stage60[20], stage60[21]},
      {stage62[0], stage62[1], stage62[2], stage62[3], stage62[4], stage62[5]},
      {stage64[0], stage63[65], stage62[66], stage61[73], stage60[90]}
   );
   gpc606_5 gpc606_5_960(
      {stage60[22], stage60[23], stage60[24], stage60[25], stage60[26], stage60[27]},
      {stage62[6], stage62[7], stage62[8], stage62[9], stage62[10], stage62[11]},
      {stage64[1], stage63[66], stage62[67], stage61[74], stage60[91]}
   );
   gpc606_5 gpc606_5_961(
      {stage60[28], stage60[29], stage60[30], stage60[31], stage60[32], stage60[33]},
      {stage62[12], stage62[13], stage62[14], stage62[15], stage62[16], stage62[17]},
      {stage64[2], stage63[67], stage62[68], stage61[75], stage60[92]}
   );
   gpc606_5 gpc606_5_962(
      {stage60[34], stage60[35], stage60[36], stage60[37], stage60[38], stage60[39]},
      {stage62[18], stage62[19], stage62[20], stage62[21], stage62[22], stage62[23]},
      {stage64[3], stage63[68], stage62[69], stage61[76], stage60[93]}
   );
   gpc606_5 gpc606_5_963(
      {stage60[40], stage60[41], stage60[42], stage60[43], stage60[44], stage60[45]},
      {stage62[24], stage62[25], stage62[26], stage62[27], stage62[28], stage62[29]},
      {stage64[4], stage63[69], stage62[70], stage61[77], stage60[94]}
   );
   gpc606_5 gpc606_5_964(
      {stage60[46], stage60[47], stage60[48], stage60[49], stage60[50], stage60[51]},
      {stage62[30], stage62[31], stage62[32], stage62[33], stage62[34], stage62[35]},
      {stage64[5], stage63[70], stage62[71], stage61[78], stage60[95]}
   );
   gpc606_5 gpc606_5_965(
      {stage60[52], stage60[53], stage60[54], stage60[55], stage60[56], stage60[57]},
      {stage62[36], stage62[37], stage62[38], stage62[39], stage62[40], stage62[41]},
      {stage64[6], stage63[71], stage62[72], stage61[79], stage60[96]}
   );
   gpc606_5 gpc606_5_966(
      {stage60[58], stage60[59], stage60[60], stage60[61], stage60[62], stage60[63]},
      {stage62[42], stage62[43], stage62[44], stage62[45], stage62[46], stage62[47]},
      {stage64[7], stage63[72], stage62[73], stage61[80], stage60[97]}
   );
   gpc1_1 gpc1_1_967(
      {stage61[6]},
      {stage61[81]}
   );
   gpc1_1 gpc1_1_968(
      {stage61[7]},
      {stage61[82]}
   );
   gpc1_1 gpc1_1_969(
      {stage61[8]},
      {stage61[83]}
   );
   gpc1_1 gpc1_1_970(
      {stage61[9]},
      {stage61[84]}
   );
   gpc1_1 gpc1_1_971(
      {stage61[10]},
      {stage61[85]}
   );
   gpc1_1 gpc1_1_972(
      {stage61[11]},
      {stage61[86]}
   );
   gpc1_1 gpc1_1_973(
      {stage61[12]},
      {stage61[87]}
   );
   gpc1_1 gpc1_1_974(
      {stage61[13]},
      {stage61[88]}
   );
   gpc1_1 gpc1_1_975(
      {stage61[14]},
      {stage61[89]}
   );
   gpc1_1 gpc1_1_976(
      {stage61[15]},
      {stage61[90]}
   );
   gpc1_1 gpc1_1_977(
      {stage61[16]},
      {stage61[91]}
   );
   gpc1_1 gpc1_1_978(
      {stage61[17]},
      {stage61[92]}
   );
   gpc1_1 gpc1_1_979(
      {stage61[18]},
      {stage61[93]}
   );
   gpc1_1 gpc1_1_980(
      {stage61[19]},
      {stage61[94]}
   );
   gpc1_1 gpc1_1_981(
      {stage61[20]},
      {stage61[95]}
   );
   gpc606_5 gpc606_5_982(
      {stage61[21], stage61[22], stage61[23], stage61[24], stage61[25], stage61[26]},
      {stage63[0], stage63[1], stage63[2], stage63[3], stage63[4], stage63[5]},
      {stage65[0], stage64[8], stage63[73], stage62[74], stage61[96]}
   );
   gpc606_5 gpc606_5_983(
      {stage61[27], stage61[28], stage61[29], stage61[30], stage61[31], stage61[32]},
      {stage63[6], stage63[7], stage63[8], stage63[9], stage63[10], stage63[11]},
      {stage65[1], stage64[9], stage63[74], stage62[75], stage61[97]}
   );
   gpc606_5 gpc606_5_984(
      {stage61[33], stage61[34], stage61[35], stage61[36], stage61[37], stage61[38]},
      {stage63[12], stage63[13], stage63[14], stage63[15], stage63[16], stage63[17]},
      {stage65[2], stage64[10], stage63[75], stage62[76], stage61[98]}
   );
   gpc615_5 gpc615_5_985(
      {stage61[39], stage61[40], stage61[41], stage61[42], stage61[43]},
      {stage62[48]},
      {stage63[18], stage63[19], stage63[20], stage63[21], stage63[22], stage63[23]},
      {stage65[3], stage64[11], stage63[76], stage62[77], stage61[99]}
   );
   gpc615_5 gpc615_5_986(
      {stage61[44], stage61[45], stage61[46], stage61[47], stage61[48]},
      {stage62[49]},
      {stage63[24], stage63[25], stage63[26], stage63[27], stage63[28], stage63[29]},
      {stage65[4], stage64[12], stage63[77], stage62[78], stage61[100]}
   );
   gpc615_5 gpc615_5_987(
      {stage61[49], stage61[50], stage61[51], stage61[52], stage61[53]},
      {stage62[50]},
      {stage63[30], stage63[31], stage63[32], stage63[33], stage63[34], stage63[35]},
      {stage65[5], stage64[13], stage63[78], stage62[79], stage61[101]}
   );
   gpc615_5 gpc615_5_988(
      {stage61[54], stage61[55], stage61[56], stage61[57], stage61[58]},
      {stage62[51]},
      {stage63[36], stage63[37], stage63[38], stage63[39], stage63[40], stage63[41]},
      {stage65[6], stage64[14], stage63[79], stage62[80], stage61[102]}
   );
   gpc615_5 gpc615_5_989(
      {stage61[59], stage61[60], stage61[61], stage61[62], stage61[63]},
      {stage62[52]},
      {stage63[42], stage63[43], stage63[44], stage63[45], stage63[46], stage63[47]},
      {stage65[7], stage64[15], stage63[80], stage62[81], stage61[103]}
   );
   gpc1_1 gpc1_1_990(
      {stage62[53]},
      {stage62[82]}
   );
   gpc1_1 gpc1_1_991(
      {stage62[54]},
      {stage62[83]}
   );
   gpc1_1 gpc1_1_992(
      {stage62[55]},
      {stage62[84]}
   );
   gpc1_1 gpc1_1_993(
      {stage62[56]},
      {stage62[85]}
   );
   gpc1_1 gpc1_1_994(
      {stage62[57]},
      {stage62[86]}
   );
   gpc1_1 gpc1_1_995(
      {stage62[58]},
      {stage62[87]}
   );
   gpc1_1 gpc1_1_996(
      {stage62[59]},
      {stage62[88]}
   );
   gpc1_1 gpc1_1_997(
      {stage62[60]},
      {stage62[89]}
   );
   gpc1_1 gpc1_1_998(
      {stage62[61]},
      {stage62[90]}
   );
   gpc1_1 gpc1_1_999(
      {stage62[62]},
      {stage62[91]}
   );
   gpc1_1 gpc1_1_1000(
      {stage62[63]},
      {stage62[92]}
   );
   gpc1_1 gpc1_1_1001(
      {stage63[48]},
      {stage63[81]}
   );
   gpc1_1 gpc1_1_1002(
      {stage63[49]},
      {stage63[82]}
   );
   gpc1_1 gpc1_1_1003(
      {stage63[50]},
      {stage63[83]}
   );
   gpc1_1 gpc1_1_1004(
      {stage63[51]},
      {stage63[84]}
   );
   gpc1_1 gpc1_1_1005(
      {stage63[52]},
      {stage63[85]}
   );
   gpc1_1 gpc1_1_1006(
      {stage63[53]},
      {stage63[86]}
   );
   gpc1_1 gpc1_1_1007(
      {stage63[54]},
      {stage63[87]}
   );
   gpc1_1 gpc1_1_1008(
      {stage63[55]},
      {stage63[88]}
   );
   gpc1_1 gpc1_1_1009(
      {stage63[56]},
      {stage63[89]}
   );
   gpc1_1 gpc1_1_1010(
      {stage63[57]},
      {stage63[90]}
   );
   gpc1_1 gpc1_1_1011(
      {stage63[58]},
      {stage63[91]}
   );
   gpc1_1 gpc1_1_1012(
      {stage63[59]},
      {stage63[92]}
   );
   gpc1_1 gpc1_1_1013(
      {stage63[60]},
      {stage63[93]}
   );
   gpc1_1 gpc1_1_1014(
      {stage63[61]},
      {stage63[94]}
   );
   gpc1_1 gpc1_1_1015(
      {stage63[62]},
      {stage63[95]}
   );
   gpc1_1 gpc1_1_1016(
      {stage63[63]},
      {stage63[96]}
   );
   gpc1_1 gpc1_1_1017(
      {stage00[64]},
      {stage00[80]}
   );
   gpc1_1 gpc1_1_1018(
      {stage00[65]},
      {stage00[81]}
   );
   gpc1_1 gpc1_1_1019(
      {stage00[66]},
      {stage00[82]}
   );
   gpc1_1 gpc1_1_1020(
      {stage00[67]},
      {stage00[83]}
   );
   gpc606_5 gpc606_5_1021(
      {stage00[68], stage00[69], stage00[70], stage00[71], stage00[72], stage00[73]},
      {stage02[64], stage02[65], stage02[66], stage02[67], stage02[68], stage02[69]},
      {stage04[93], stage03[121], stage02[86], stage01[110], stage00[84]}
   );
   gpc606_5 gpc606_5_1022(
      {stage00[74], stage00[75], stage00[76], stage00[77], stage00[78], stage00[79]},
      {stage02[70], stage02[71], stage02[72], stage02[73], stage02[74], stage02[75]},
      {stage04[94], stage03[122], stage02[87], stage01[111], stage00[85]}
   );
   gpc1_1 gpc1_1_1023(
      {stage01[64]},
      {stage01[112]}
   );
   gpc1_1 gpc1_1_1024(
      {stage01[65]},
      {stage01[113]}
   );
   gpc1_1 gpc1_1_1025(
      {stage01[66]},
      {stage01[114]}
   );
   gpc1_1 gpc1_1_1026(
      {stage01[67]},
      {stage01[115]}
   );
   gpc606_5 gpc606_5_1027(
      {stage01[68], stage01[69], stage01[70], stage01[71], stage01[72], stage01[73]},
      {stage03[64], stage03[65], stage03[66], stage03[67], stage03[68], stage03[69]},
      {stage05[90], stage04[95], stage03[123], stage02[88], stage01[116]}
   );
   gpc606_5 gpc606_5_1028(
      {stage01[74], stage01[75], stage01[76], stage01[77], stage01[78], stage01[79]},
      {stage03[70], stage03[71], stage03[72], stage03[73], stage03[74], stage03[75]},
      {stage05[91], stage04[96], stage03[124], stage02[89], stage01[117]}
   );
   gpc606_5 gpc606_5_1029(
      {stage01[80], stage01[81], stage01[82], stage01[83], stage01[84], stage01[85]},
      {stage03[76], stage03[77], stage03[78], stage03[79], stage03[80], stage03[81]},
      {stage05[92], stage04[97], stage03[125], stage02[90], stage01[118]}
   );
   gpc606_5 gpc606_5_1030(
      {stage01[86], stage01[87], stage01[88], stage01[89], stage01[90], stage01[91]},
      {stage03[82], stage03[83], stage03[84], stage03[85], stage03[86], stage03[87]},
      {stage05[93], stage04[98], stage03[126], stage02[91], stage01[119]}
   );
   gpc606_5 gpc606_5_1031(
      {stage01[92], stage01[93], stage01[94], stage01[95], stage01[96], stage01[97]},
      {stage03[88], stage03[89], stage03[90], stage03[91], stage03[92], stage03[93]},
      {stage05[94], stage04[99], stage03[127], stage02[92], stage01[120]}
   );
   gpc606_5 gpc606_5_1032(
      {stage01[98], stage01[99], stage01[100], stage01[101], stage01[102], stage01[103]},
      {stage03[94], stage03[95], stage03[96], stage03[97], stage03[98], stage03[99]},
      {stage05[95], stage04[100], stage03[128], stage02[93], stage01[121]}
   );
   gpc606_5 gpc606_5_1033(
      {stage01[104], stage01[105], stage01[106], stage01[107], stage01[108], stage01[109]},
      {stage03[100], stage03[101], stage03[102], stage03[103], stage03[104], stage03[105]},
      {stage05[96], stage04[101], stage03[129], stage02[94], stage01[122]}
   );
   gpc1_1 gpc1_1_1034(
      {stage02[76]},
      {stage02[95]}
   );
   gpc1_1 gpc1_1_1035(
      {stage02[77]},
      {stage02[96]}
   );
   gpc1_1 gpc1_1_1036(
      {stage02[78]},
      {stage02[97]}
   );
   gpc1_1 gpc1_1_1037(
      {stage02[79]},
      {stage02[98]}
   );
   gpc1_1 gpc1_1_1038(
      {stage02[80]},
      {stage02[99]}
   );
   gpc1_1 gpc1_1_1039(
      {stage02[81]},
      {stage02[100]}
   );
   gpc1_1 gpc1_1_1040(
      {stage02[82]},
      {stage02[101]}
   );
   gpc1_1 gpc1_1_1041(
      {stage02[83]},
      {stage02[102]}
   );
   gpc1_1 gpc1_1_1042(
      {stage02[84]},
      {stage02[103]}
   );
   gpc1_1 gpc1_1_1043(
      {stage02[85]},
      {stage02[104]}
   );
   gpc615_5 gpc615_5_1044(
      {stage03[106], stage03[107], stage03[108], stage03[109], stage03[110]},
      {stage04[64]},
      {stage05[64], stage05[65], stage05[66], stage05[67], stage05[68], stage05[69]},
      {stage07[97], stage06[90], stage05[97], stage04[102], stage03[130]}
   );
   gpc615_5 gpc615_5_1045(
      {stage03[111], stage03[112], stage03[113], stage03[114], stage03[115]},
      {stage04[65]},
      {stage05[70], stage05[71], stage05[72], stage05[73], stage05[74], stage05[75]},
      {stage07[98], stage06[91], stage05[98], stage04[103], stage03[131]}
   );
   gpc615_5 gpc615_5_1046(
      {stage03[116], stage03[117], stage03[118], stage03[119], stage03[120]},
      {stage04[66]},
      {stage05[76], stage05[77], stage05[78], stage05[79], stage05[80], stage05[81]},
      {stage07[99], stage06[92], stage05[99], stage04[104], stage03[132]}
   );
   gpc1_1 gpc1_1_1047(
      {stage04[67]},
      {stage04[105]}
   );
   gpc1_1 gpc1_1_1048(
      {stage04[68]},
      {stage04[106]}
   );
   gpc1_1 gpc1_1_1049(
      {stage04[69]},
      {stage04[107]}
   );
   gpc606_5 gpc606_5_1050(
      {stage04[70], stage04[71], stage04[72], stage04[73], stage04[74], stage04[75]},
      {stage06[64], stage06[65], stage06[66], stage06[67], stage06[68], stage06[69]},
      {stage08[102], stage07[100], stage06[93], stage05[100], stage04[108]}
   );
   gpc606_5 gpc606_5_1051(
      {stage04[76], stage04[77], stage04[78], stage04[79], stage04[80], stage04[81]},
      {stage06[70], stage06[71], stage06[72], stage06[73], stage06[74], stage06[75]},
      {stage08[103], stage07[101], stage06[94], stage05[101], stage04[109]}
   );
   gpc606_5 gpc606_5_1052(
      {stage04[82], stage04[83], stage04[84], stage04[85], stage04[86], stage04[87]},
      {stage06[76], stage06[77], stage06[78], stage06[79], stage06[80], stage06[81]},
      {stage08[104], stage07[102], stage06[95], stage05[102], stage04[110]}
   );
   gpc615_5 gpc615_5_1053(
      {stage04[88], stage04[89], stage04[90], stage04[91], stage04[92]},
      {stage05[82]},
      {stage06[82], stage06[83], stage06[84], stage06[85], stage06[86], stage06[87]},
      {stage08[105], stage07[103], stage06[96], stage05[103], stage04[111]}
   );
   gpc1_1 gpc1_1_1054(
      {stage05[83]},
      {stage05[104]}
   );
   gpc1_1 gpc1_1_1055(
      {stage05[84]},
      {stage05[105]}
   );
   gpc1_1 gpc1_1_1056(
      {stage05[85]},
      {stage05[106]}
   );
   gpc1_1 gpc1_1_1057(
      {stage05[86]},
      {stage05[107]}
   );
   gpc1_1 gpc1_1_1058(
      {stage05[87]},
      {stage05[108]}
   );
   gpc1_1 gpc1_1_1059(
      {stage05[88]},
      {stage05[109]}
   );
   gpc1_1 gpc1_1_1060(
      {stage05[89]},
      {stage05[110]}
   );
   gpc1_1 gpc1_1_1061(
      {stage06[88]},
      {stage06[97]}
   );
   gpc1_1 gpc1_1_1062(
      {stage06[89]},
      {stage06[98]}
   );
   gpc615_5 gpc615_5_1063(
      {stage07[64], stage07[65], stage07[66], stage07[67], stage07[68]},
      {stage08[64]},
      {stage09[64], stage09[65], stage09[66], stage09[67], stage09[68], stage09[69]},
      {stage11[93], stage10[110], stage09[123], stage08[106], stage07[104]}
   );
   gpc615_5 gpc615_5_1064(
      {stage07[69], stage07[70], stage07[71], stage07[72], stage07[73]},
      {stage08[65]},
      {stage09[70], stage09[71], stage09[72], stage09[73], stage09[74], stage09[75]},
      {stage11[94], stage10[111], stage09[124], stage08[107], stage07[105]}
   );
   gpc615_5 gpc615_5_1065(
      {stage07[74], stage07[75], stage07[76], stage07[77], stage07[78]},
      {stage08[66]},
      {stage09[76], stage09[77], stage09[78], stage09[79], stage09[80], stage09[81]},
      {stage11[95], stage10[112], stage09[125], stage08[108], stage07[106]}
   );
   gpc615_5 gpc615_5_1066(
      {stage07[79], stage07[80], stage07[81], stage07[82], stage07[83]},
      {stage08[67]},
      {stage09[82], stage09[83], stage09[84], stage09[85], stage09[86], stage09[87]},
      {stage11[96], stage10[113], stage09[126], stage08[109], stage07[107]}
   );
   gpc615_5 gpc615_5_1067(
      {stage07[84], stage07[85], stage07[86], stage07[87], stage07[88]},
      {stage08[68]},
      {stage09[88], stage09[89], stage09[90], stage09[91], stage09[92], stage09[93]},
      {stage11[97], stage10[114], stage09[127], stage08[110], stage07[108]}
   );
   gpc615_5 gpc615_5_1068(
      {stage07[89], stage07[90], stage07[91], stage07[92], stage07[93]},
      {stage08[69]},
      {stage09[94], stage09[95], stage09[96], stage09[97], stage09[98], stage09[99]},
      {stage11[98], stage10[115], stage09[128], stage08[111], stage07[109]}
   );
   gpc615_5 gpc615_5_1069(
      {stage07[94], stage07[95], stage07[96], 1'h0, 1'h0},
      {stage08[70]},
      {stage09[100], stage09[101], stage09[102], stage09[103], stage09[104], stage09[105]},
      {stage11[99], stage10[116], stage09[129], stage08[112], stage07[110]}
   );
   gpc1_1 gpc1_1_1070(
      {stage08[71]},
      {stage08[113]}
   );
   gpc606_5 gpc606_5_1071(
      {stage08[72], stage08[73], stage08[74], stage08[75], stage08[76], stage08[77]},
      {stage10[64], stage10[65], stage10[66], stage10[67], stage10[68], stage10[69]},
      {stage12[110], stage11[100], stage10[117], stage09[130], stage08[114]}
   );
   gpc606_5 gpc606_5_1072(
      {stage08[78], stage08[79], stage08[80], stage08[81], stage08[82], stage08[83]},
      {stage10[70], stage10[71], stage10[72], stage10[73], stage10[74], stage10[75]},
      {stage12[111], stage11[101], stage10[118], stage09[131], stage08[115]}
   );
   gpc606_5 gpc606_5_1073(
      {stage08[84], stage08[85], stage08[86], stage08[87], stage08[88], stage08[89]},
      {stage10[76], stage10[77], stage10[78], stage10[79], stage10[80], stage10[81]},
      {stage12[112], stage11[102], stage10[119], stage09[132], stage08[116]}
   );
   gpc606_5 gpc606_5_1074(
      {stage08[90], stage08[91], stage08[92], stage08[93], stage08[94], stage08[95]},
      {stage10[82], stage10[83], stage10[84], stage10[85], stage10[86], stage10[87]},
      {stage12[113], stage11[103], stage10[120], stage09[133], stage08[117]}
   );
   gpc606_5 gpc606_5_1075(
      {stage08[96], stage08[97], stage08[98], stage08[99], stage08[100], stage08[101]},
      {stage10[88], stage10[89], stage10[90], stage10[91], stage10[92], stage10[93]},
      {stage12[114], stage11[104], stage10[121], stage09[134], stage08[118]}
   );
   gpc1_1 gpc1_1_1076(
      {stage09[106]},
      {stage09[135]}
   );
   gpc1_1 gpc1_1_1077(
      {stage09[107]},
      {stage09[136]}
   );
   gpc1_1 gpc1_1_1078(
      {stage09[108]},
      {stage09[137]}
   );
   gpc1_1 gpc1_1_1079(
      {stage09[109]},
      {stage09[138]}
   );
   gpc1_1 gpc1_1_1080(
      {stage09[110]},
      {stage09[139]}
   );
   gpc1_1 gpc1_1_1081(
      {stage09[111]},
      {stage09[140]}
   );
   gpc1_1 gpc1_1_1082(
      {stage09[112]},
      {stage09[141]}
   );
   gpc1_1 gpc1_1_1083(
      {stage09[113]},
      {stage09[142]}
   );
   gpc1_1 gpc1_1_1084(
      {stage09[114]},
      {stage09[143]}
   );
   gpc1_1 gpc1_1_1085(
      {stage09[115]},
      {stage09[144]}
   );
   gpc1_1 gpc1_1_1086(
      {stage09[116]},
      {stage09[145]}
   );
   gpc1_1 gpc1_1_1087(
      {stage09[117]},
      {stage09[146]}
   );
   gpc1_1 gpc1_1_1088(
      {stage09[118]},
      {stage09[147]}
   );
   gpc1_1 gpc1_1_1089(
      {stage09[119]},
      {stage09[148]}
   );
   gpc1_1 gpc1_1_1090(
      {stage09[120]},
      {stage09[149]}
   );
   gpc1_1 gpc1_1_1091(
      {stage09[121]},
      {stage09[150]}
   );
   gpc1_1 gpc1_1_1092(
      {stage09[122]},
      {stage09[151]}
   );
   gpc1_1 gpc1_1_1093(
      {stage10[94]},
      {stage10[122]}
   );
   gpc1_1 gpc1_1_1094(
      {stage10[95]},
      {stage10[123]}
   );
   gpc1_1 gpc1_1_1095(
      {stage10[96]},
      {stage10[124]}
   );
   gpc1_1 gpc1_1_1096(
      {stage10[97]},
      {stage10[125]}
   );
   gpc1_1 gpc1_1_1097(
      {stage10[98]},
      {stage10[126]}
   );
   gpc1_1 gpc1_1_1098(
      {stage10[99]},
      {stage10[127]}
   );
   gpc615_5 gpc615_5_1099(
      {stage10[100], stage10[101], stage10[102], stage10[103], stage10[104]},
      {stage11[64]},
      {stage12[64], stage12[65], stage12[66], stage12[67], stage12[68], stage12[69]},
      {stage14[94], stage13[90], stage12[115], stage11[105], stage10[128]}
   );
   gpc615_5 gpc615_5_1100(
      {stage10[105], stage10[106], stage10[107], stage10[108], stage10[109]},
      {stage11[65]},
      {stage12[70], stage12[71], stage12[72], stage12[73], stage12[74], stage12[75]},
      {stage14[95], stage13[91], stage12[116], stage11[106], stage10[129]}
   );
   gpc1_1 gpc1_1_1101(
      {stage11[66]},
      {stage11[107]}
   );
   gpc1_1 gpc1_1_1102(
      {stage11[67]},
      {stage11[108]}
   );
   gpc1_1 gpc1_1_1103(
      {stage11[68]},
      {stage11[109]}
   );
   gpc1_1 gpc1_1_1104(
      {stage11[69]},
      {stage11[110]}
   );
   gpc1_1 gpc1_1_1105(
      {stage11[70]},
      {stage11[111]}
   );
   gpc1_1 gpc1_1_1106(
      {stage11[71]},
      {stage11[112]}
   );
   gpc1_1 gpc1_1_1107(
      {stage11[72]},
      {stage11[113]}
   );
   gpc1_1 gpc1_1_1108(
      {stage11[73]},
      {stage11[114]}
   );
   gpc1_1 gpc1_1_1109(
      {stage11[74]},
      {stage11[115]}
   );
   gpc1_1 gpc1_1_1110(
      {stage11[75]},
      {stage11[116]}
   );
   gpc1_1 gpc1_1_1111(
      {stage11[76]},
      {stage11[117]}
   );
   gpc1_1 gpc1_1_1112(
      {stage11[77]},
      {stage11[118]}
   );
   gpc1_1 gpc1_1_1113(
      {stage11[78]},
      {stage11[119]}
   );
   gpc1_1 gpc1_1_1114(
      {stage11[79]},
      {stage11[120]}
   );
   gpc1_1 gpc1_1_1115(
      {stage11[80]},
      {stage11[121]}
   );
   gpc1_1 gpc1_1_1116(
      {stage11[81]},
      {stage11[122]}
   );
   gpc1_1 gpc1_1_1117(
      {stage11[82]},
      {stage11[123]}
   );
   gpc1_1 gpc1_1_1118(
      {stage11[83]},
      {stage11[124]}
   );
   gpc1_1 gpc1_1_1119(
      {stage11[84]},
      {stage11[125]}
   );
   gpc1_1 gpc1_1_1120(
      {stage11[85]},
      {stage11[126]}
   );
   gpc1_1 gpc1_1_1121(
      {stage11[86]},
      {stage11[127]}
   );
   gpc1_1 gpc1_1_1122(
      {stage11[87]},
      {stage11[128]}
   );
   gpc1_1 gpc1_1_1123(
      {stage11[88]},
      {stage11[129]}
   );
   gpc1_1 gpc1_1_1124(
      {stage11[89]},
      {stage11[130]}
   );
   gpc1_1 gpc1_1_1125(
      {stage11[90]},
      {stage11[131]}
   );
   gpc1_1 gpc1_1_1126(
      {stage11[91]},
      {stage11[132]}
   );
   gpc1_1 gpc1_1_1127(
      {stage11[92]},
      {stage11[133]}
   );
   gpc1_1 gpc1_1_1128(
      {stage12[76]},
      {stage12[117]}
   );
   gpc1_1 gpc1_1_1129(
      {stage12[77]},
      {stage12[118]}
   );
   gpc1_1 gpc1_1_1130(
      {stage12[78]},
      {stage12[119]}
   );
   gpc1_1 gpc1_1_1131(
      {stage12[79]},
      {stage12[120]}
   );
   gpc1_1 gpc1_1_1132(
      {stage12[80]},
      {stage12[121]}
   );
   gpc1_1 gpc1_1_1133(
      {stage12[81]},
      {stage12[122]}
   );
   gpc1_1 gpc1_1_1134(
      {stage12[82]},
      {stage12[123]}
   );
   gpc1_1 gpc1_1_1135(
      {stage12[83]},
      {stage12[124]}
   );
   gpc1_1 gpc1_1_1136(
      {stage12[84]},
      {stage12[125]}
   );
   gpc1_1 gpc1_1_1137(
      {stage12[85]},
      {stage12[126]}
   );
   gpc606_5 gpc606_5_1138(
      {stage12[86], stage12[87], stage12[88], stage12[89], stage12[90], stage12[91]},
      {stage14[64], stage14[65], stage14[66], stage14[67], stage14[68], stage14[69]},
      {stage16[90], stage15[124], stage14[96], stage13[92], stage12[127]}
   );
   gpc606_5 gpc606_5_1139(
      {stage12[92], stage12[93], stage12[94], stage12[95], stage12[96], stage12[97]},
      {stage14[70], stage14[71], stage14[72], stage14[73], stage14[74], stage14[75]},
      {stage16[91], stage15[125], stage14[97], stage13[93], stage12[128]}
   );
   gpc606_5 gpc606_5_1140(
      {stage12[98], stage12[99], stage12[100], stage12[101], stage12[102], stage12[103]},
      {stage14[76], stage14[77], stage14[78], stage14[79], stage14[80], stage14[81]},
      {stage16[92], stage15[126], stage14[98], stage13[94], stage12[129]}
   );
   gpc606_5 gpc606_5_1141(
      {stage12[104], stage12[105], stage12[106], stage12[107], stage12[108], stage12[109]},
      {stage14[82], stage14[83], stage14[84], stage14[85], stage14[86], stage14[87]},
      {stage16[93], stage15[127], stage14[99], stage13[95], stage12[130]}
   );
   gpc1_1 gpc1_1_1142(
      {stage13[64]},
      {stage13[96]}
   );
   gpc1_1 gpc1_1_1143(
      {stage13[65]},
      {stage13[97]}
   );
   gpc1_1 gpc1_1_1144(
      {stage13[66]},
      {stage13[98]}
   );
   gpc1_1 gpc1_1_1145(
      {stage13[67]},
      {stage13[99]}
   );
   gpc1_1 gpc1_1_1146(
      {stage13[68]},
      {stage13[100]}
   );
   gpc1_1 gpc1_1_1147(
      {stage13[69]},
      {stage13[101]}
   );
   gpc1_1 gpc1_1_1148(
      {stage13[70]},
      {stage13[102]}
   );
   gpc1_1 gpc1_1_1149(
      {stage13[71]},
      {stage13[103]}
   );
   gpc606_5 gpc606_5_1150(
      {stage13[72], stage13[73], stage13[74], stage13[75], stage13[76], stage13[77]},
      {stage15[64], stage15[65], stage15[66], stage15[67], stage15[68], stage15[69]},
      {stage17[104], stage16[94], stage15[128], stage14[100], stage13[104]}
   );
   gpc606_5 gpc606_5_1151(
      {stage13[78], stage13[79], stage13[80], stage13[81], stage13[82], stage13[83]},
      {stage15[70], stage15[71], stage15[72], stage15[73], stage15[74], stage15[75]},
      {stage17[105], stage16[95], stage15[129], stage14[101], stage13[105]}
   );
   gpc606_5 gpc606_5_1152(
      {stage13[84], stage13[85], stage13[86], stage13[87], stage13[88], stage13[89]},
      {stage15[76], stage15[77], stage15[78], stage15[79], stage15[80], stage15[81]},
      {stage17[106], stage16[96], stage15[130], stage14[102], stage13[106]}
   );
   gpc1_1 gpc1_1_1153(
      {stage14[88]},
      {stage14[103]}
   );
   gpc615_5 gpc615_5_1154(
      {stage14[89], stage14[90], stage14[91], stage14[92], stage14[93]},
      {stage15[82]},
      {stage16[64], stage16[65], stage16[66], stage16[67], stage16[68], stage16[69]},
      {stage18[85], stage17[107], stage16[97], stage15[131], stage14[104]}
   );
   gpc1_1 gpc1_1_1155(
      {stage15[83]},
      {stage15[132]}
   );
   gpc1_1 gpc1_1_1156(
      {stage15[84]},
      {stage15[133]}
   );
   gpc1_1 gpc1_1_1157(
      {stage15[85]},
      {stage15[134]}
   );
   gpc1_1 gpc1_1_1158(
      {stage15[86]},
      {stage15[135]}
   );
   gpc1_1 gpc1_1_1159(
      {stage15[87]},
      {stage15[136]}
   );
   gpc1_1 gpc1_1_1160(
      {stage15[88]},
      {stage15[137]}
   );
   gpc2135_5 gpc2135_5_1161(
      {stage15[89], stage15[90], stage15[91], stage15[92], stage15[93]},
      {stage16[70], stage16[71], stage16[72]},
      {stage17[64]},
      {stage18[64], stage18[65]},
      {stage19[99], stage18[86], stage17[108], stage16[98], stage15[138]}
   );
   gpc2135_5 gpc2135_5_1162(
      {stage15[94], stage15[95], stage15[96], stage15[97], stage15[98]},
      {stage16[73], stage16[74], stage16[75]},
      {stage17[65]},
      {stage18[66], stage18[67]},
      {stage19[100], stage18[87], stage17[109], stage16[99], stage15[139]}
   );
   gpc2135_5 gpc2135_5_1163(
      {stage15[99], stage15[100], stage15[101], stage15[102], stage15[103]},
      {stage16[76], stage16[77], stage16[78]},
      {stage17[66]},
      {stage18[68], stage18[69]},
      {stage19[101], stage18[88], stage17[110], stage16[100], stage15[140]}
   );
   gpc2135_5 gpc2135_5_1164(
      {stage15[104], stage15[105], stage15[106], stage15[107], stage15[108]},
      {stage16[79], stage16[80], stage16[81]},
      {stage17[67]},
      {stage18[70], stage18[71]},
      {stage19[102], stage18[89], stage17[111], stage16[101], stage15[141]}
   );
   gpc2135_5 gpc2135_5_1165(
      {stage15[109], stage15[110], stage15[111], stage15[112], stage15[113]},
      {stage16[82], stage16[83], stage16[84]},
      {stage17[68]},
      {stage18[72], stage18[73]},
      {stage19[103], stage18[90], stage17[112], stage16[102], stage15[142]}
   );
   gpc2135_5 gpc2135_5_1166(
      {stage15[114], stage15[115], stage15[116], stage15[117], stage15[118]},
      {stage16[85], stage16[86], stage16[87]},
      {stage17[69]},
      {stage18[74], stage18[75]},
      {stage19[104], stage18[91], stage17[113], stage16[103], stage15[143]}
   );
   gpc2135_5 gpc2135_5_1167(
      {stage15[119], stage15[120], stage15[121], stage15[122], stage15[123]},
      {stage16[88], stage16[89], 1'h0},
      {stage17[70]},
      {stage18[76], stage18[77]},
      {stage19[105], stage18[92], stage17[114], stage16[104], stage15[144]}
   );
   gpc1_1 gpc1_1_1168(
      {stage17[71]},
      {stage17[115]}
   );
   gpc1_1 gpc1_1_1169(
      {stage17[72]},
      {stage17[116]}
   );
   gpc1_1 gpc1_1_1170(
      {stage17[73]},
      {stage17[117]}
   );
   gpc1_1 gpc1_1_1171(
      {stage17[74]},
      {stage17[118]}
   );
   gpc1_1 gpc1_1_1172(
      {stage17[75]},
      {stage17[119]}
   );
   gpc1_1 gpc1_1_1173(
      {stage17[76]},
      {stage17[120]}
   );
   gpc1_1 gpc1_1_1174(
      {stage17[77]},
      {stage17[121]}
   );
   gpc1_1 gpc1_1_1175(
      {stage17[78]},
      {stage17[122]}
   );
   gpc1_1 gpc1_1_1176(
      {stage17[79]},
      {stage17[123]}
   );
   gpc1_1 gpc1_1_1177(
      {stage17[80]},
      {stage17[124]}
   );
   gpc1_1 gpc1_1_1178(
      {stage17[81]},
      {stage17[125]}
   );
   gpc1_1 gpc1_1_1179(
      {stage17[82]},
      {stage17[126]}
   );
   gpc1_1 gpc1_1_1180(
      {stage17[83]},
      {stage17[127]}
   );
   gpc1_1 gpc1_1_1181(
      {stage17[84]},
      {stage17[128]}
   );
   gpc1_1 gpc1_1_1182(
      {stage17[85]},
      {stage17[129]}
   );
   gpc1_1 gpc1_1_1183(
      {stage17[86]},
      {stage17[130]}
   );
   gpc1_1 gpc1_1_1184(
      {stage17[87]},
      {stage17[131]}
   );
   gpc1_1 gpc1_1_1185(
      {stage17[88]},
      {stage17[132]}
   );
   gpc1_1 gpc1_1_1186(
      {stage17[89]},
      {stage17[133]}
   );
   gpc1_1 gpc1_1_1187(
      {stage17[90]},
      {stage17[134]}
   );
   gpc1_1 gpc1_1_1188(
      {stage17[91]},
      {stage17[135]}
   );
   gpc606_5 gpc606_5_1189(
      {stage17[92], stage17[93], stage17[94], stage17[95], stage17[96], stage17[97]},
      {stage19[64], stage19[65], stage19[66], stage19[67], stage19[68], stage19[69]},
      {stage21[91], stage20[106], stage19[106], stage18[93], stage17[136]}
   );
   gpc606_5 gpc606_5_1190(
      {stage17[98], stage17[99], stage17[100], stage17[101], stage17[102], stage17[103]},
      {stage19[70], stage19[71], stage19[72], stage19[73], stage19[74], stage19[75]},
      {stage21[92], stage20[107], stage19[107], stage18[94], stage17[137]}
   );
   gpc1_1 gpc1_1_1191(
      {stage18[78]},
      {stage18[95]}
   );
   gpc1_1 gpc1_1_1192(
      {stage18[79]},
      {stage18[96]}
   );
   gpc1_1 gpc1_1_1193(
      {stage18[80]},
      {stage18[97]}
   );
   gpc1_1 gpc1_1_1194(
      {stage18[81]},
      {stage18[98]}
   );
   gpc1_1 gpc1_1_1195(
      {stage18[82]},
      {stage18[99]}
   );
   gpc1_1 gpc1_1_1196(
      {stage18[83]},
      {stage18[100]}
   );
   gpc1_1 gpc1_1_1197(
      {stage18[84]},
      {stage18[101]}
   );
   gpc1_1 gpc1_1_1198(
      {stage19[76]},
      {stage19[108]}
   );
   gpc1_1 gpc1_1_1199(
      {stage19[77]},
      {stage19[109]}
   );
   gpc1_1 gpc1_1_1200(
      {stage19[78]},
      {stage19[110]}
   );
   gpc615_5 gpc615_5_1201(
      {stage19[79], stage19[80], stage19[81], stage19[82], stage19[83]},
      {stage20[64]},
      {stage21[64], stage21[65], stage21[66], stage21[67], stage21[68], stage21[69]},
      {stage23[95], stage22[99], stage21[93], stage20[108], stage19[111]}
   );
   gpc615_5 gpc615_5_1202(
      {stage19[84], stage19[85], stage19[86], stage19[87], stage19[88]},
      {stage20[65]},
      {stage21[70], stage21[71], stage21[72], stage21[73], stage21[74], stage21[75]},
      {stage23[96], stage22[100], stage21[94], stage20[109], stage19[112]}
   );
   gpc615_5 gpc615_5_1203(
      {stage19[89], stage19[90], stage19[91], stage19[92], stage19[93]},
      {stage20[66]},
      {stage21[76], stage21[77], stage21[78], stage21[79], stage21[80], stage21[81]},
      {stage23[97], stage22[101], stage21[95], stage20[110], stage19[113]}
   );
   gpc615_5 gpc615_5_1204(
      {stage19[94], stage19[95], stage19[96], stage19[97], stage19[98]},
      {stage20[67]},
      {stage21[82], stage21[83], stage21[84], stage21[85], stage21[86], stage21[87]},
      {stage23[98], stage22[102], stage21[96], stage20[111], stage19[114]}
   );
   gpc1_1 gpc1_1_1205(
      {stage20[68]},
      {stage20[112]}
   );
   gpc1_1 gpc1_1_1206(
      {stage20[69]},
      {stage20[113]}
   );
   gpc1_1 gpc1_1_1207(
      {stage20[70]},
      {stage20[114]}
   );
   gpc1_1 gpc1_1_1208(
      {stage20[71]},
      {stage20[115]}
   );
   gpc1_1 gpc1_1_1209(
      {stage20[72]},
      {stage20[116]}
   );
   gpc1_1 gpc1_1_1210(
      {stage20[73]},
      {stage20[117]}
   );
   gpc1_1 gpc1_1_1211(
      {stage20[74]},
      {stage20[118]}
   );
   gpc1_1 gpc1_1_1212(
      {stage20[75]},
      {stage20[119]}
   );
   gpc606_5 gpc606_5_1213(
      {stage20[76], stage20[77], stage20[78], stage20[79], stage20[80], stage20[81]},
      {stage22[64], stage22[65], stage22[66], stage22[67], stage22[68], stage22[69]},
      {stage24[98], stage23[99], stage22[103], stage21[97], stage20[120]}
   );
   gpc606_5 gpc606_5_1214(
      {stage20[82], stage20[83], stage20[84], stage20[85], stage20[86], stage20[87]},
      {stage22[70], stage22[71], stage22[72], stage22[73], stage22[74], stage22[75]},
      {stage24[99], stage23[100], stage22[104], stage21[98], stage20[121]}
   );
   gpc606_5 gpc606_5_1215(
      {stage20[88], stage20[89], stage20[90], stage20[91], stage20[92], stage20[93]},
      {stage22[76], stage22[77], stage22[78], stage22[79], stage22[80], stage22[81]},
      {stage24[100], stage23[101], stage22[105], stage21[99], stage20[122]}
   );
   gpc606_5 gpc606_5_1216(
      {stage20[94], stage20[95], stage20[96], stage20[97], stage20[98], stage20[99]},
      {stage22[82], stage22[83], stage22[84], stage22[85], stage22[86], stage22[87]},
      {stage24[101], stage23[102], stage22[106], stage21[100], stage20[123]}
   );
   gpc606_5 gpc606_5_1217(
      {stage20[100], stage20[101], stage20[102], stage20[103], stage20[104], stage20[105]},
      {stage22[88], stage22[89], stage22[90], stage22[91], stage22[92], stage22[93]},
      {stage24[102], stage23[103], stage22[107], stage21[101], stage20[124]}
   );
   gpc1_1 gpc1_1_1218(
      {stage21[88]},
      {stage21[102]}
   );
   gpc1_1 gpc1_1_1219(
      {stage21[89]},
      {stage21[103]}
   );
   gpc1_1 gpc1_1_1220(
      {stage21[90]},
      {stage21[104]}
   );
   gpc615_5 gpc615_5_1221(
      {stage22[94], stage22[95], stage22[96], stage22[97], stage22[98]},
      {stage23[64]},
      {stage24[64], stage24[65], stage24[66], stage24[67], stage24[68], stage24[69]},
      {stage26[87], stage25[98], stage24[103], stage23[104], stage22[108]}
   );
   gpc1_1 gpc1_1_1222(
      {stage23[65]},
      {stage23[105]}
   );
   gpc1_1 gpc1_1_1223(
      {stage23[66]},
      {stage23[106]}
   );
   gpc1_1 gpc1_1_1224(
      {stage23[67]},
      {stage23[107]}
   );
   gpc1_1 gpc1_1_1225(
      {stage23[68]},
      {stage23[108]}
   );
   gpc1_1 gpc1_1_1226(
      {stage23[69]},
      {stage23[109]}
   );
   gpc1_1 gpc1_1_1227(
      {stage23[70]},
      {stage23[110]}
   );
   gpc1_1 gpc1_1_1228(
      {stage23[71]},
      {stage23[111]}
   );
   gpc1_1 gpc1_1_1229(
      {stage23[72]},
      {stage23[112]}
   );
   gpc1_1 gpc1_1_1230(
      {stage23[73]},
      {stage23[113]}
   );
   gpc1_1 gpc1_1_1231(
      {stage23[74]},
      {stage23[114]}
   );
   gpc615_5 gpc615_5_1232(
      {stage23[75], stage23[76], stage23[77], stage23[78], stage23[79]},
      {stage24[70]},
      {stage25[64], stage25[65], stage25[66], stage25[67], stage25[68], stage25[69]},
      {stage27[104], stage26[88], stage25[99], stage24[104], stage23[115]}
   );
   gpc615_5 gpc615_5_1233(
      {stage23[80], stage23[81], stage23[82], stage23[83], stage23[84]},
      {stage24[71]},
      {stage25[70], stage25[71], stage25[72], stage25[73], stage25[74], stage25[75]},
      {stage27[105], stage26[89], stage25[100], stage24[105], stage23[116]}
   );
   gpc615_5 gpc615_5_1234(
      {stage23[85], stage23[86], stage23[87], stage23[88], stage23[89]},
      {stage24[72]},
      {stage25[76], stage25[77], stage25[78], stage25[79], stage25[80], stage25[81]},
      {stage27[106], stage26[90], stage25[101], stage24[106], stage23[117]}
   );
   gpc615_5 gpc615_5_1235(
      {stage23[90], stage23[91], stage23[92], stage23[93], stage23[94]},
      {stage24[73]},
      {stage25[82], stage25[83], stage25[84], stage25[85], stage25[86], stage25[87]},
      {stage27[107], stage26[91], stage25[102], stage24[107], stage23[118]}
   );
   gpc606_5 gpc606_5_1236(
      {stage24[74], stage24[75], stage24[76], stage24[77], stage24[78], stage24[79]},
      {stage26[64], stage26[65], stage26[66], stage26[67], stage26[68], stage26[69]},
      {stage28[90], stage27[108], stage26[92], stage25[103], stage24[108]}
   );
   gpc606_5 gpc606_5_1237(
      {stage24[80], stage24[81], stage24[82], stage24[83], stage24[84], stage24[85]},
      {stage26[70], stage26[71], stage26[72], stage26[73], stage26[74], stage26[75]},
      {stage28[91], stage27[109], stage26[93], stage25[104], stage24[109]}
   );
   gpc606_5 gpc606_5_1238(
      {stage24[86], stage24[87], stage24[88], stage24[89], stage24[90], stage24[91]},
      {stage26[76], stage26[77], stage26[78], stage26[79], stage26[80], stage26[81]},
      {stage28[92], stage27[110], stage26[94], stage25[105], stage24[110]}
   );
   gpc606_5 gpc606_5_1239(
      {stage24[92], stage24[93], stage24[94], stage24[95], stage24[96], stage24[97]},
      {stage26[82], stage26[83], stage26[84], stage26[85], stage26[86], 1'h0},
      {stage28[93], stage27[111], stage26[95], stage25[106], stage24[111]}
   );
   gpc1_1 gpc1_1_1240(
      {stage25[88]},
      {stage25[107]}
   );
   gpc1_1 gpc1_1_1241(
      {stage25[89]},
      {stage25[108]}
   );
   gpc1_1 gpc1_1_1242(
      {stage25[90]},
      {stage25[109]}
   );
   gpc1_1 gpc1_1_1243(
      {stage25[91]},
      {stage25[110]}
   );
   gpc1_1 gpc1_1_1244(
      {stage25[92]},
      {stage25[111]}
   );
   gpc1_1 gpc1_1_1245(
      {stage25[93]},
      {stage25[112]}
   );
   gpc1_1 gpc1_1_1246(
      {stage25[94]},
      {stage25[113]}
   );
   gpc1_1 gpc1_1_1247(
      {stage25[95]},
      {stage25[114]}
   );
   gpc1_1 gpc1_1_1248(
      {stage25[96]},
      {stage25[115]}
   );
   gpc1_1 gpc1_1_1249(
      {stage25[97]},
      {stage25[116]}
   );
   gpc1_1 gpc1_1_1250(
      {stage27[64]},
      {stage27[112]}
   );
   gpc1_1 gpc1_1_1251(
      {stage27[65]},
      {stage27[113]}
   );
   gpc1_1 gpc1_1_1252(
      {stage27[66]},
      {stage27[114]}
   );
   gpc1_1 gpc1_1_1253(
      {stage27[67]},
      {stage27[115]}
   );
   gpc1_1 gpc1_1_1254(
      {stage27[68]},
      {stage27[116]}
   );
   gpc1_1 gpc1_1_1255(
      {stage27[69]},
      {stage27[117]}
   );
   gpc1_1 gpc1_1_1256(
      {stage27[70]},
      {stage27[118]}
   );
   gpc1_1 gpc1_1_1257(
      {stage27[71]},
      {stage27[119]}
   );
   gpc1_1 gpc1_1_1258(
      {stage27[72]},
      {stage27[120]}
   );
   gpc1_1 gpc1_1_1259(
      {stage27[73]},
      {stage27[121]}
   );
   gpc606_5 gpc606_5_1260(
      {stage27[74], stage27[75], stage27[76], stage27[77], stage27[78], stage27[79]},
      {stage29[64], stage29[65], stage29[66], stage29[67], stage29[68], stage29[69]},
      {stage31[91], stage30[94], stage29[94], stage28[94], stage27[122]}
   );
   gpc606_5 gpc606_5_1261(
      {stage27[80], stage27[81], stage27[82], stage27[83], stage27[84], stage27[85]},
      {stage29[70], stage29[71], stage29[72], stage29[73], stage29[74], stage29[75]},
      {stage31[92], stage30[95], stage29[95], stage28[95], stage27[123]}
   );
   gpc606_5 gpc606_5_1262(
      {stage27[86], stage27[87], stage27[88], stage27[89], stage27[90], stage27[91]},
      {stage29[76], stage29[77], stage29[78], stage29[79], stage29[80], stage29[81]},
      {stage31[93], stage30[96], stage29[96], stage28[96], stage27[124]}
   );
   gpc606_5 gpc606_5_1263(
      {stage27[92], stage27[93], stage27[94], stage27[95], stage27[96], stage27[97]},
      {stage29[82], stage29[83], stage29[84], stage29[85], stage29[86], stage29[87]},
      {stage31[94], stage30[97], stage29[97], stage28[97], stage27[125]}
   );
   gpc606_5 gpc606_5_1264(
      {stage27[98], stage27[99], stage27[100], stage27[101], stage27[102], stage27[103]},
      {stage29[88], stage29[89], stage29[90], stage29[91], stage29[92], stage29[93]},
      {stage31[95], stage30[98], stage29[98], stage28[98], stage27[126]}
   );
   gpc1_1 gpc1_1_1265(
      {stage28[64]},
      {stage28[99]}
   );
   gpc1_1 gpc1_1_1266(
      {stage28[65]},
      {stage28[100]}
   );
   gpc1_1 gpc1_1_1267(
      {stage28[66]},
      {stage28[101]}
   );
   gpc1_1 gpc1_1_1268(
      {stage28[67]},
      {stage28[102]}
   );
   gpc1_1 gpc1_1_1269(
      {stage28[68]},
      {stage28[103]}
   );
   gpc1_1 gpc1_1_1270(
      {stage28[69]},
      {stage28[104]}
   );
   gpc1_1 gpc1_1_1271(
      {stage28[70]},
      {stage28[105]}
   );
   gpc1_1 gpc1_1_1272(
      {stage28[71]},
      {stage28[106]}
   );
   gpc1_1 gpc1_1_1273(
      {stage28[72]},
      {stage28[107]}
   );
   gpc1_1 gpc1_1_1274(
      {stage28[73]},
      {stage28[108]}
   );
   gpc1_1 gpc1_1_1275(
      {stage28[74]},
      {stage28[109]}
   );
   gpc1_1 gpc1_1_1276(
      {stage28[75]},
      {stage28[110]}
   );
   gpc1_1 gpc1_1_1277(
      {stage28[76]},
      {stage28[111]}
   );
   gpc1_1 gpc1_1_1278(
      {stage28[77]},
      {stage28[112]}
   );
   gpc1_1 gpc1_1_1279(
      {stage28[78]},
      {stage28[113]}
   );
   gpc1_1 gpc1_1_1280(
      {stage28[79]},
      {stage28[114]}
   );
   gpc1_1 gpc1_1_1281(
      {stage28[80]},
      {stage28[115]}
   );
   gpc1_1 gpc1_1_1282(
      {stage28[81]},
      {stage28[116]}
   );
   gpc1_1 gpc1_1_1283(
      {stage28[82]},
      {stage28[117]}
   );
   gpc1_1 gpc1_1_1284(
      {stage28[83]},
      {stage28[118]}
   );
   gpc1_1 gpc1_1_1285(
      {stage28[84]},
      {stage28[119]}
   );
   gpc1_1 gpc1_1_1286(
      {stage28[85]},
      {stage28[120]}
   );
   gpc1_1 gpc1_1_1287(
      {stage28[86]},
      {stage28[121]}
   );
   gpc1_1 gpc1_1_1288(
      {stage28[87]},
      {stage28[122]}
   );
   gpc1_1 gpc1_1_1289(
      {stage28[88]},
      {stage28[123]}
   );
   gpc1_1 gpc1_1_1290(
      {stage28[89]},
      {stage28[124]}
   );
   gpc1_1 gpc1_1_1291(
      {stage30[64]},
      {stage30[99]}
   );
   gpc1_1 gpc1_1_1292(
      {stage30[65]},
      {stage30[100]}
   );
   gpc1_1 gpc1_1_1293(
      {stage30[66]},
      {stage30[101]}
   );
   gpc1_1 gpc1_1_1294(
      {stage30[67]},
      {stage30[102]}
   );
   gpc1_1 gpc1_1_1295(
      {stage30[68]},
      {stage30[103]}
   );
   gpc1_1 gpc1_1_1296(
      {stage30[69]},
      {stage30[104]}
   );
   gpc1_1 gpc1_1_1297(
      {stage30[70]},
      {stage30[105]}
   );
   gpc1_1 gpc1_1_1298(
      {stage30[71]},
      {stage30[106]}
   );
   gpc1_1 gpc1_1_1299(
      {stage30[72]},
      {stage30[107]}
   );
   gpc1_1 gpc1_1_1300(
      {stage30[73]},
      {stage30[108]}
   );
   gpc1_1 gpc1_1_1301(
      {stage30[74]},
      {stage30[109]}
   );
   gpc1_1 gpc1_1_1302(
      {stage30[75]},
      {stage30[110]}
   );
   gpc1_1 gpc1_1_1303(
      {stage30[76]},
      {stage30[111]}
   );
   gpc1_1 gpc1_1_1304(
      {stage30[77]},
      {stage30[112]}
   );
   gpc1_1 gpc1_1_1305(
      {stage30[78]},
      {stage30[113]}
   );
   gpc1_1 gpc1_1_1306(
      {stage30[79]},
      {stage30[114]}
   );
   gpc1_1 gpc1_1_1307(
      {stage30[80]},
      {stage30[115]}
   );
   gpc1_1 gpc1_1_1308(
      {stage30[81]},
      {stage30[116]}
   );
   gpc623_5 gpc623_5_1309(
      {stage30[82], stage30[83], stage30[84]},
      {stage31[64], stage31[65]},
      {stage32[64], stage32[65], stage32[66], stage32[67], stage32[68], stage32[69]},
      {stage34[88], stage33[90], stage32[97], stage31[96], stage30[117]}
   );
   gpc623_5 gpc623_5_1310(
      {stage30[85], stage30[86], stage30[87]},
      {stage31[66], stage31[67]},
      {stage32[70], stage32[71], stage32[72], stage32[73], stage32[74], stage32[75]},
      {stage34[89], stage33[91], stage32[98], stage31[97], stage30[118]}
   );
   gpc623_5 gpc623_5_1311(
      {stage30[88], stage30[89], stage30[90]},
      {stage31[68], stage31[69]},
      {stage32[76], stage32[77], stage32[78], stage32[79], stage32[80], stage32[81]},
      {stage34[90], stage33[92], stage32[99], stage31[98], stage30[119]}
   );
   gpc623_5 gpc623_5_1312(
      {stage30[91], stage30[92], stage30[93]},
      {stage31[70], stage31[71]},
      {stage32[82], stage32[83], stage32[84], stage32[85], stage32[86], stage32[87]},
      {stage34[91], stage33[93], stage32[100], stage31[99], stage30[120]}
   );
   gpc1_1 gpc1_1_1313(
      {stage31[72]},
      {stage31[100]}
   );
   gpc1_1 gpc1_1_1314(
      {stage31[73]},
      {stage31[101]}
   );
   gpc1_1 gpc1_1_1315(
      {stage31[74]},
      {stage31[102]}
   );
   gpc1_1 gpc1_1_1316(
      {stage31[75]},
      {stage31[103]}
   );
   gpc615_5 gpc615_5_1317(
      {stage31[76], stage31[77], stage31[78], stage31[79], stage31[80]},
      {stage32[88]},
      {stage33[64], stage33[65], stage33[66], stage33[67], stage33[68], stage33[69]},
      {stage35[91], stage34[92], stage33[94], stage32[101], stage31[104]}
   );
   gpc615_5 gpc615_5_1318(
      {stage31[81], stage31[82], stage31[83], stage31[84], stage31[85]},
      {stage32[89]},
      {stage33[70], stage33[71], stage33[72], stage33[73], stage33[74], stage33[75]},
      {stage35[92], stage34[93], stage33[95], stage32[102], stage31[105]}
   );
   gpc615_5 gpc615_5_1319(
      {stage31[86], stage31[87], stage31[88], stage31[89], stage31[90]},
      {stage32[90]},
      {stage33[76], stage33[77], stage33[78], stage33[79], stage33[80], stage33[81]},
      {stage35[93], stage34[94], stage33[96], stage32[103], stage31[106]}
   );
   gpc606_5 gpc606_5_1320(
      {stage32[91], stage32[92], stage32[93], stage32[94], stage32[95], stage32[96]},
      {stage34[64], stage34[65], stage34[66], stage34[67], stage34[68], stage34[69]},
      {stage36[107], stage35[94], stage34[95], stage33[97], stage32[104]}
   );
   gpc1_1 gpc1_1_1321(
      {stage33[82]},
      {stage33[98]}
   );
   gpc1_1 gpc1_1_1322(
      {stage33[83]},
      {stage33[99]}
   );
   gpc1_1 gpc1_1_1323(
      {stage33[84]},
      {stage33[100]}
   );
   gpc1_1 gpc1_1_1324(
      {stage33[85]},
      {stage33[101]}
   );
   gpc1_1 gpc1_1_1325(
      {stage33[86]},
      {stage33[102]}
   );
   gpc1_1 gpc1_1_1326(
      {stage33[87]},
      {stage33[103]}
   );
   gpc1_1 gpc1_1_1327(
      {stage33[88]},
      {stage33[104]}
   );
   gpc1_1 gpc1_1_1328(
      {stage33[89]},
      {stage33[105]}
   );
   gpc1_1 gpc1_1_1329(
      {stage34[70]},
      {stage34[96]}
   );
   gpc1_1 gpc1_1_1330(
      {stage34[71]},
      {stage34[97]}
   );
   gpc1_1 gpc1_1_1331(
      {stage34[72]},
      {stage34[98]}
   );
   gpc615_5 gpc615_5_1332(
      {stage34[73], stage34[74], stage34[75], stage34[76], stage34[77]},
      {stage35[64]},
      {stage36[64], stage36[65], stage36[66], stage36[67], stage36[68], stage36[69]},
      {stage38[88], stage37[96], stage36[108], stage35[95], stage34[99]}
   );
   gpc615_5 gpc615_5_1333(
      {stage34[78], stage34[79], stage34[80], stage34[81], stage34[82]},
      {stage35[65]},
      {stage36[70], stage36[71], stage36[72], stage36[73], stage36[74], stage36[75]},
      {stage38[89], stage37[97], stage36[109], stage35[96], stage34[100]}
   );
   gpc615_5 gpc615_5_1334(
      {stage34[83], stage34[84], stage34[85], stage34[86], stage34[87]},
      {stage35[66]},
      {stage36[76], stage36[77], stage36[78], stage36[79], stage36[80], stage36[81]},
      {stage38[90], stage37[98], stage36[110], stage35[97], stage34[101]}
   );
   gpc1_1 gpc1_1_1335(
      {stage35[67]},
      {stage35[98]}
   );
   gpc1_1 gpc1_1_1336(
      {stage35[68]},
      {stage35[99]}
   );
   gpc1_1 gpc1_1_1337(
      {stage35[69]},
      {stage35[100]}
   );
   gpc1_1 gpc1_1_1338(
      {stage35[70]},
      {stage35[101]}
   );
   gpc615_5 gpc615_5_1339(
      {stage35[71], stage35[72], stage35[73], stage35[74], stage35[75]},
      {stage36[82]},
      {stage37[64], stage37[65], stage37[66], stage37[67], stage37[68], stage37[69]},
      {stage39[92], stage38[91], stage37[99], stage36[111], stage35[102]}
   );
   gpc615_5 gpc615_5_1340(
      {stage35[76], stage35[77], stage35[78], stage35[79], stage35[80]},
      {stage36[83]},
      {stage37[70], stage37[71], stage37[72], stage37[73], stage37[74], stage37[75]},
      {stage39[93], stage38[92], stage37[100], stage36[112], stage35[103]}
   );
   gpc615_5 gpc615_5_1341(
      {stage35[81], stage35[82], stage35[83], stage35[84], stage35[85]},
      {stage36[84]},
      {stage37[76], stage37[77], stage37[78], stage37[79], stage37[80], stage37[81]},
      {stage39[94], stage38[93], stage37[101], stage36[113], stage35[104]}
   );
   gpc615_5 gpc615_5_1342(
      {stage35[86], stage35[87], stage35[88], stage35[89], stage35[90]},
      {stage36[85]},
      {stage37[82], stage37[83], stage37[84], stage37[85], stage37[86], stage37[87]},
      {stage39[95], stage38[94], stage37[102], stage36[114], stage35[105]}
   );
   gpc1_1 gpc1_1_1343(
      {stage36[86]},
      {stage36[115]}
   );
   gpc1_1 gpc1_1_1344(
      {stage36[87]},
      {stage36[116]}
   );
   gpc1_1 gpc1_1_1345(
      {stage36[88]},
      {stage36[117]}
   );
   gpc606_5 gpc606_5_1346(
      {stage36[89], stage36[90], stage36[91], stage36[92], stage36[93], stage36[94]},
      {stage38[64], stage38[65], stage38[66], stage38[67], stage38[68], stage38[69]},
      {stage40[101], stage39[96], stage38[95], stage37[103], stage36[118]}
   );
   gpc606_5 gpc606_5_1347(
      {stage36[95], stage36[96], stage36[97], stage36[98], stage36[99], stage36[100]},
      {stage38[70], stage38[71], stage38[72], stage38[73], stage38[74], stage38[75]},
      {stage40[102], stage39[97], stage38[96], stage37[104], stage36[119]}
   );
   gpc606_5 gpc606_5_1348(
      {stage36[101], stage36[102], stage36[103], stage36[104], stage36[105], stage36[106]},
      {stage38[76], stage38[77], stage38[78], stage38[79], stage38[80], stage38[81]},
      {stage40[103], stage39[98], stage38[97], stage37[105], stage36[120]}
   );
   gpc1_1 gpc1_1_1349(
      {stage37[88]},
      {stage37[106]}
   );
   gpc1_1 gpc1_1_1350(
      {stage37[89]},
      {stage37[107]}
   );
   gpc1406_5 gpc1406_5_1351(
      {stage37[90], stage37[91], stage37[92], stage37[93], stage37[94], stage37[95]},
      {stage39[64], stage39[65], stage39[66], stage39[67]},
      {stage40[64]},
      {stage41[110], stage40[104], stage39[99], stage38[98], stage37[108]}
   );
   gpc1_1 gpc1_1_1352(
      {stage38[82]},
      {stage38[99]}
   );
   gpc1_1 gpc1_1_1353(
      {stage38[83]},
      {stage38[100]}
   );
   gpc1_1 gpc1_1_1354(
      {stage38[84]},
      {stage38[101]}
   );
   gpc1_1 gpc1_1_1355(
      {stage38[85]},
      {stage38[102]}
   );
   gpc1_1 gpc1_1_1356(
      {stage38[86]},
      {stage38[103]}
   );
   gpc1_1 gpc1_1_1357(
      {stage38[87]},
      {stage38[104]}
   );
   gpc606_5 gpc606_5_1358(
      {stage39[68], stage39[69], stage39[70], stage39[71], stage39[72], stage39[73]},
      {stage41[64], stage41[65], stage41[66], stage41[67], stage41[68], stage41[69]},
      {stage43[99], stage42[106], stage41[111], stage40[105], stage39[100]}
   );
   gpc606_5 gpc606_5_1359(
      {stage39[74], stage39[75], stage39[76], stage39[77], stage39[78], stage39[79]},
      {stage41[70], stage41[71], stage41[72], stage41[73], stage41[74], stage41[75]},
      {stage43[100], stage42[107], stage41[112], stage40[106], stage39[101]}
   );
   gpc606_5 gpc606_5_1360(
      {stage39[80], stage39[81], stage39[82], stage39[83], stage39[84], stage39[85]},
      {stage41[76], stage41[77], stage41[78], stage41[79], stage41[80], stage41[81]},
      {stage43[101], stage42[108], stage41[113], stage40[107], stage39[102]}
   );
   gpc606_5 gpc606_5_1361(
      {stage39[86], stage39[87], stage39[88], stage39[89], stage39[90], stage39[91]},
      {stage41[82], stage41[83], stage41[84], stage41[85], stage41[86], stage41[87]},
      {stage43[102], stage42[109], stage41[114], stage40[108], stage39[103]}
   );
   gpc1_1 gpc1_1_1362(
      {stage40[65]},
      {stage40[109]}
   );
   gpc1_1 gpc1_1_1363(
      {stage40[66]},
      {stage40[110]}
   );
   gpc1_1 gpc1_1_1364(
      {stage40[67]},
      {stage40[111]}
   );
   gpc1_1 gpc1_1_1365(
      {stage40[68]},
      {stage40[112]}
   );
   gpc1_1 gpc1_1_1366(
      {stage40[69]},
      {stage40[113]}
   );
   gpc1_1 gpc1_1_1367(
      {stage40[70]},
      {stage40[114]}
   );
   gpc606_5 gpc606_5_1368(
      {stage40[71], stage40[72], stage40[73], stage40[74], stage40[75], stage40[76]},
      {stage42[64], stage42[65], stage42[66], stage42[67], stage42[68], stage42[69]},
      {stage44[85], stage43[103], stage42[110], stage41[115], stage40[115]}
   );
   gpc606_5 gpc606_5_1369(
      {stage40[77], stage40[78], stage40[79], stage40[80], stage40[81], stage40[82]},
      {stage42[70], stage42[71], stage42[72], stage42[73], stage42[74], stage42[75]},
      {stage44[86], stage43[104], stage42[111], stage41[116], stage40[116]}
   );
   gpc606_5 gpc606_5_1370(
      {stage40[83], stage40[84], stage40[85], stage40[86], stage40[87], stage40[88]},
      {stage42[76], stage42[77], stage42[78], stage42[79], stage42[80], stage42[81]},
      {stage44[87], stage43[105], stage42[112], stage41[117], stage40[117]}
   );
   gpc606_5 gpc606_5_1371(
      {stage40[89], stage40[90], stage40[91], stage40[92], stage40[93], stage40[94]},
      {stage42[82], stage42[83], stage42[84], stage42[85], stage42[86], stage42[87]},
      {stage44[88], stage43[106], stage42[113], stage41[118], stage40[118]}
   );
   gpc606_5 gpc606_5_1372(
      {stage40[95], stage40[96], stage40[97], stage40[98], stage40[99], stage40[100]},
      {stage42[88], stage42[89], stage42[90], stage42[91], stage42[92], stage42[93]},
      {stage44[89], stage43[107], stage42[114], stage41[119], stage40[119]}
   );
   gpc1_1 gpc1_1_1373(
      {stage41[88]},
      {stage41[120]}
   );
   gpc1_1 gpc1_1_1374(
      {stage41[89]},
      {stage41[121]}
   );
   gpc1_1 gpc1_1_1375(
      {stage41[90]},
      {stage41[122]}
   );
   gpc1_1 gpc1_1_1376(
      {stage41[91]},
      {stage41[123]}
   );
   gpc606_5 gpc606_5_1377(
      {stage41[92], stage41[93], stage41[94], stage41[95], stage41[96], stage41[97]},
      {stage43[64], stage43[65], stage43[66], stage43[67], stage43[68], stage43[69]},
      {stage45[93], stage44[90], stage43[108], stage42[115], stage41[124]}
   );
   gpc606_5 gpc606_5_1378(
      {stage41[98], stage41[99], stage41[100], stage41[101], stage41[102], stage41[103]},
      {stage43[70], stage43[71], stage43[72], stage43[73], stage43[74], stage43[75]},
      {stage45[94], stage44[91], stage43[109], stage42[116], stage41[125]}
   );
   gpc606_5 gpc606_5_1379(
      {stage41[104], stage41[105], stage41[106], stage41[107], stage41[108], stage41[109]},
      {stage43[76], stage43[77], stage43[78], stage43[79], stage43[80], stage43[81]},
      {stage45[95], stage44[92], stage43[110], stage42[117], stage41[126]}
   );
   gpc1_1 gpc1_1_1380(
      {stage42[94]},
      {stage42[118]}
   );
   gpc1_1 gpc1_1_1381(
      {stage42[95]},
      {stage42[119]}
   );
   gpc1_1 gpc1_1_1382(
      {stage42[96]},
      {stage42[120]}
   );
   gpc1_1 gpc1_1_1383(
      {stage42[97]},
      {stage42[121]}
   );
   gpc1_1 gpc1_1_1384(
      {stage42[98]},
      {stage42[122]}
   );
   gpc1_1 gpc1_1_1385(
      {stage42[99]},
      {stage42[123]}
   );
   gpc1_1 gpc1_1_1386(
      {stage42[100]},
      {stage42[124]}
   );
   gpc1_1 gpc1_1_1387(
      {stage42[101]},
      {stage42[125]}
   );
   gpc1_1 gpc1_1_1388(
      {stage42[102]},
      {stage42[126]}
   );
   gpc1_1 gpc1_1_1389(
      {stage42[103]},
      {stage42[127]}
   );
   gpc1_1 gpc1_1_1390(
      {stage42[104]},
      {stage42[128]}
   );
   gpc1_1 gpc1_1_1391(
      {stage42[105]},
      {stage42[129]}
   );
   gpc1_1 gpc1_1_1392(
      {stage43[82]},
      {stage43[111]}
   );
   gpc1_1 gpc1_1_1393(
      {stage43[83]},
      {stage43[112]}
   );
   gpc1_1 gpc1_1_1394(
      {stage43[84]},
      {stage43[113]}
   );
   gpc1_1 gpc1_1_1395(
      {stage43[85]},
      {stage43[114]}
   );
   gpc1_1 gpc1_1_1396(
      {stage43[86]},
      {stage43[115]}
   );
   gpc1_1 gpc1_1_1397(
      {stage43[87]},
      {stage43[116]}
   );
   gpc1_1 gpc1_1_1398(
      {stage43[88]},
      {stage43[117]}
   );
   gpc1_1 gpc1_1_1399(
      {stage43[89]},
      {stage43[118]}
   );
   gpc1_1 gpc1_1_1400(
      {stage43[90]},
      {stage43[119]}
   );
   gpc1_1 gpc1_1_1401(
      {stage43[91]},
      {stage43[120]}
   );
   gpc1_1 gpc1_1_1402(
      {stage43[92]},
      {stage43[121]}
   );
   gpc1_1 gpc1_1_1403(
      {stage43[93]},
      {stage43[122]}
   );
   gpc1_1 gpc1_1_1404(
      {stage43[94]},
      {stage43[123]}
   );
   gpc1_1 gpc1_1_1405(
      {stage43[95]},
      {stage43[124]}
   );
   gpc1_1 gpc1_1_1406(
      {stage43[96]},
      {stage43[125]}
   );
   gpc1_1 gpc1_1_1407(
      {stage43[97]},
      {stage43[126]}
   );
   gpc1_1 gpc1_1_1408(
      {stage43[98]},
      {stage43[127]}
   );
   gpc1_1 gpc1_1_1409(
      {stage44[64]},
      {stage44[93]}
   );
   gpc1_1 gpc1_1_1410(
      {stage44[65]},
      {stage44[94]}
   );
   gpc1_1 gpc1_1_1411(
      {stage44[66]},
      {stage44[95]}
   );
   gpc1_1 gpc1_1_1412(
      {stage44[67]},
      {stage44[96]}
   );
   gpc1_1 gpc1_1_1413(
      {stage44[68]},
      {stage44[97]}
   );
   gpc1_1 gpc1_1_1414(
      {stage44[69]},
      {stage44[98]}
   );
   gpc1_1 gpc1_1_1415(
      {stage44[70]},
      {stage44[99]}
   );
   gpc1_1 gpc1_1_1416(
      {stage44[71]},
      {stage44[100]}
   );
   gpc1_1 gpc1_1_1417(
      {stage44[72]},
      {stage44[101]}
   );
   gpc1_1 gpc1_1_1418(
      {stage44[73]},
      {stage44[102]}
   );
   gpc1_1 gpc1_1_1419(
      {stage44[74]},
      {stage44[103]}
   );
   gpc1_1 gpc1_1_1420(
      {stage44[75]},
      {stage44[104]}
   );
   gpc1_1 gpc1_1_1421(
      {stage44[76]},
      {stage44[105]}
   );
   gpc1_1 gpc1_1_1422(
      {stage44[77]},
      {stage44[106]}
   );
   gpc1_1 gpc1_1_1423(
      {stage44[78]},
      {stage44[107]}
   );
   gpc606_5 gpc606_5_1424(
      {stage44[79], stage44[80], stage44[81], stage44[82], stage44[83], stage44[84]},
      {stage46[64], stage46[65], stage46[66], stage46[67], stage46[68], stage46[69]},
      {stage48[101], stage47[91], stage46[106], stage45[96], stage44[108]}
   );
   gpc1_1 gpc1_1_1425(
      {stage45[64]},
      {stage45[97]}
   );
   gpc1_1 gpc1_1_1426(
      {stage45[65]},
      {stage45[98]}
   );
   gpc1_1 gpc1_1_1427(
      {stage45[66]},
      {stage45[99]}
   );
   gpc1_1 gpc1_1_1428(
      {stage45[67]},
      {stage45[100]}
   );
   gpc1_1 gpc1_1_1429(
      {stage45[68]},
      {stage45[101]}
   );
   gpc1_1 gpc1_1_1430(
      {stage45[69]},
      {stage45[102]}
   );
   gpc1_1 gpc1_1_1431(
      {stage45[70]},
      {stage45[103]}
   );
   gpc1_1 gpc1_1_1432(
      {stage45[71]},
      {stage45[104]}
   );
   gpc1_1 gpc1_1_1433(
      {stage45[72]},
      {stage45[105]}
   );
   gpc1_1 gpc1_1_1434(
      {stage45[73]},
      {stage45[106]}
   );
   gpc1_1 gpc1_1_1435(
      {stage45[74]},
      {stage45[107]}
   );
   gpc1_1 gpc1_1_1436(
      {stage45[75]},
      {stage45[108]}
   );
   gpc1_1 gpc1_1_1437(
      {stage45[76]},
      {stage45[109]}
   );
   gpc1_1 gpc1_1_1438(
      {stage45[77]},
      {stage45[110]}
   );
   gpc1_1 gpc1_1_1439(
      {stage45[78]},
      {stage45[111]}
   );
   gpc1_1 gpc1_1_1440(
      {stage45[79]},
      {stage45[112]}
   );
   gpc1_1 gpc1_1_1441(
      {stage45[80]},
      {stage45[113]}
   );
   gpc1_1 gpc1_1_1442(
      {stage45[81]},
      {stage45[114]}
   );
   gpc1_1 gpc1_1_1443(
      {stage45[82]},
      {stage45[115]}
   );
   gpc1_1 gpc1_1_1444(
      {stage45[83]},
      {stage45[116]}
   );
   gpc1_1 gpc1_1_1445(
      {stage45[84]},
      {stage45[117]}
   );
   gpc1_1 gpc1_1_1446(
      {stage45[85]},
      {stage45[118]}
   );
   gpc1_1 gpc1_1_1447(
      {stage45[86]},
      {stage45[119]}
   );
   gpc1_1 gpc1_1_1448(
      {stage45[87]},
      {stage45[120]}
   );
   gpc615_5 gpc615_5_1449(
      {stage45[88], stage45[89], stage45[90], stage45[91], stage45[92]},
      {stage46[70]},
      {stage47[64], stage47[65], stage47[66], stage47[67], stage47[68], stage47[69]},
      {stage49[89], stage48[102], stage47[92], stage46[107], stage45[121]}
   );
   gpc1_1 gpc1_1_1450(
      {stage46[71]},
      {stage46[108]}
   );
   gpc1_1 gpc1_1_1451(
      {stage46[72]},
      {stage46[109]}
   );
   gpc1_1 gpc1_1_1452(
      {stage46[73]},
      {stage46[110]}
   );
   gpc1_1 gpc1_1_1453(
      {stage46[74]},
      {stage46[111]}
   );
   gpc7_3 gpc7_3_1454(
      {stage46[75], stage46[76], stage46[77], stage46[78], stage46[79], stage46[80], stage46[81]},
      {stage48[103], stage47[93], stage46[112]}
   );
   gpc7_3 gpc7_3_1455(
      {stage46[82], stage46[83], stage46[84], stage46[85], stage46[86], stage46[87], stage46[88]},
      {stage48[104], stage47[94], stage46[113]}
   );
   gpc7_3 gpc7_3_1456(
      {stage46[89], stage46[90], stage46[91], stage46[92], stage46[93], stage46[94], stage46[95]},
      {stage48[105], stage47[95], stage46[114]}
   );
   gpc615_5 gpc615_5_1457(
      {stage46[96], stage46[97], stage46[98], stage46[99], stage46[100]},
      {stage47[70]},
      {stage48[64], stage48[65], stage48[66], stage48[67], stage48[68], stage48[69]},
      {stage50[96], stage49[90], stage48[106], stage47[96], stage46[115]}
   );
   gpc615_5 gpc615_5_1458(
      {stage46[101], stage46[102], stage46[103], stage46[104], stage46[105]},
      {stage47[71]},
      {stage48[70], stage48[71], stage48[72], stage48[73], stage48[74], stage48[75]},
      {stage50[97], stage49[91], stage48[107], stage47[97], stage46[116]}
   );
   gpc1_1 gpc1_1_1459(
      {stage47[72]},
      {stage47[98]}
   );
   gpc1_1 gpc1_1_1460(
      {stage47[73]},
      {stage47[99]}
   );
   gpc1_1 gpc1_1_1461(
      {stage47[74]},
      {stage47[100]}
   );
   gpc1_1 gpc1_1_1462(
      {stage47[75]},
      {stage47[101]}
   );
   gpc1_1 gpc1_1_1463(
      {stage47[76]},
      {stage47[102]}
   );
   gpc1_1 gpc1_1_1464(
      {stage47[77]},
      {stage47[103]}
   );
   gpc1_1 gpc1_1_1465(
      {stage47[78]},
      {stage47[104]}
   );
   gpc1_1 gpc1_1_1466(
      {stage47[79]},
      {stage47[105]}
   );
   gpc1_1 gpc1_1_1467(
      {stage47[80]},
      {stage47[106]}
   );
   gpc1_1 gpc1_1_1468(
      {stage47[81]},
      {stage47[107]}
   );
   gpc1_1 gpc1_1_1469(
      {stage47[82]},
      {stage47[108]}
   );
   gpc1_1 gpc1_1_1470(
      {stage47[83]},
      {stage47[109]}
   );
   gpc1_1 gpc1_1_1471(
      {stage47[84]},
      {stage47[110]}
   );
   gpc1_1 gpc1_1_1472(
      {stage47[85]},
      {stage47[111]}
   );
   gpc1_1 gpc1_1_1473(
      {stage47[86]},
      {stage47[112]}
   );
   gpc1_1 gpc1_1_1474(
      {stage47[87]},
      {stage47[113]}
   );
   gpc1_1 gpc1_1_1475(
      {stage47[88]},
      {stage47[114]}
   );
   gpc1_1 gpc1_1_1476(
      {stage47[89]},
      {stage47[115]}
   );
   gpc1_1 gpc1_1_1477(
      {stage47[90]},
      {stage47[116]}
   );
   gpc1_1 gpc1_1_1478(
      {stage48[76]},
      {stage48[108]}
   );
   gpc606_5 gpc606_5_1479(
      {stage48[77], stage48[78], stage48[79], stage48[80], stage48[81], stage48[82]},
      {stage50[64], stage50[65], stage50[66], stage50[67], stage50[68], stage50[69]},
      {stage52[92], stage51[88], stage50[98], stage49[92], stage48[109]}
   );
   gpc606_5 gpc606_5_1480(
      {stage48[83], stage48[84], stage48[85], stage48[86], stage48[87], stage48[88]},
      {stage50[70], stage50[71], stage50[72], stage50[73], stage50[74], stage50[75]},
      {stage52[93], stage51[89], stage50[99], stage49[93], stage48[110]}
   );
   gpc606_5 gpc606_5_1481(
      {stage48[89], stage48[90], stage48[91], stage48[92], stage48[93], stage48[94]},
      {stage50[76], stage50[77], stage50[78], stage50[79], stage50[80], stage50[81]},
      {stage52[94], stage51[90], stage50[100], stage49[94], stage48[111]}
   );
   gpc606_5 gpc606_5_1482(
      {stage48[95], stage48[96], stage48[97], stage48[98], stage48[99], stage48[100]},
      {stage50[82], stage50[83], stage50[84], stage50[85], stage50[86], stage50[87]},
      {stage52[95], stage51[91], stage50[101], stage49[95], stage48[112]}
   );
   gpc1_1 gpc1_1_1483(
      {stage49[64]},
      {stage49[96]}
   );
   gpc1_1 gpc1_1_1484(
      {stage49[65]},
      {stage49[97]}
   );
   gpc1_1 gpc1_1_1485(
      {stage49[66]},
      {stage49[98]}
   );
   gpc1_1 gpc1_1_1486(
      {stage49[67]},
      {stage49[99]}
   );
   gpc1_1 gpc1_1_1487(
      {stage49[68]},
      {stage49[100]}
   );
   gpc1_1 gpc1_1_1488(
      {stage49[69]},
      {stage49[101]}
   );
   gpc1_1 gpc1_1_1489(
      {stage49[70]},
      {stage49[102]}
   );
   gpc1_1 gpc1_1_1490(
      {stage49[71]},
      {stage49[103]}
   );
   gpc1_1 gpc1_1_1491(
      {stage49[72]},
      {stage49[104]}
   );
   gpc1_1 gpc1_1_1492(
      {stage49[73]},
      {stage49[105]}
   );
   gpc1_1 gpc1_1_1493(
      {stage49[74]},
      {stage49[106]}
   );
   gpc1_1 gpc1_1_1494(
      {stage49[75]},
      {stage49[107]}
   );
   gpc1_1 gpc1_1_1495(
      {stage49[76]},
      {stage49[108]}
   );
   gpc1_1 gpc1_1_1496(
      {stage49[77]},
      {stage49[109]}
   );
   gpc1_1 gpc1_1_1497(
      {stage49[78]},
      {stage49[110]}
   );
   gpc1_1 gpc1_1_1498(
      {stage49[79]},
      {stage49[111]}
   );
   gpc1_1 gpc1_1_1499(
      {stage49[80]},
      {stage49[112]}
   );
   gpc1_1 gpc1_1_1500(
      {stage49[81]},
      {stage49[113]}
   );
   gpc1_1 gpc1_1_1501(
      {stage49[82]},
      {stage49[114]}
   );
   gpc1_1 gpc1_1_1502(
      {stage49[83]},
      {stage49[115]}
   );
   gpc615_5 gpc615_5_1503(
      {stage49[84], stage49[85], stage49[86], stage49[87], stage49[88]},
      {stage50[88]},
      {stage51[64], stage51[65], stage51[66], stage51[67], stage51[68], stage51[69]},
      {stage53[95], stage52[96], stage51[92], stage50[102], stage49[116]}
   );
   gpc1_1 gpc1_1_1504(
      {stage50[89]},
      {stage50[103]}
   );
   gpc1_1 gpc1_1_1505(
      {stage50[90]},
      {stage50[104]}
   );
   gpc1_1 gpc1_1_1506(
      {stage50[91]},
      {stage50[105]}
   );
   gpc1_1 gpc1_1_1507(
      {stage50[92]},
      {stage50[106]}
   );
   gpc1_1 gpc1_1_1508(
      {stage50[93]},
      {stage50[107]}
   );
   gpc1_1 gpc1_1_1509(
      {stage50[94]},
      {stage50[108]}
   );
   gpc1_1 gpc1_1_1510(
      {stage50[95]},
      {stage50[109]}
   );
   gpc1_1 gpc1_1_1511(
      {stage51[70]},
      {stage51[93]}
   );
   gpc1_1 gpc1_1_1512(
      {stage51[71]},
      {stage51[94]}
   );
   gpc1_1 gpc1_1_1513(
      {stage51[72]},
      {stage51[95]}
   );
   gpc1_1 gpc1_1_1514(
      {stage51[73]},
      {stage51[96]}
   );
   gpc1_1 gpc1_1_1515(
      {stage51[74]},
      {stage51[97]}
   );
   gpc1_1 gpc1_1_1516(
      {stage51[75]},
      {stage51[98]}
   );
   gpc1_1 gpc1_1_1517(
      {stage51[76]},
      {stage51[99]}
   );
   gpc1_1 gpc1_1_1518(
      {stage51[77]},
      {stage51[100]}
   );
   gpc615_5 gpc615_5_1519(
      {stage51[78], stage51[79], stage51[80], stage51[81], stage51[82]},
      {stage52[64]},
      {stage53[64], stage53[65], stage53[66], stage53[67], stage53[68], stage53[69]},
      {stage55[94], stage54[98], stage53[96], stage52[97], stage51[101]}
   );
   gpc615_5 gpc615_5_1520(
      {stage51[83], stage51[84], stage51[85], stage51[86], stage51[87]},
      {stage52[65]},
      {stage53[70], stage53[71], stage53[72], stage53[73], stage53[74], stage53[75]},
      {stage55[95], stage54[99], stage53[97], stage52[98], stage51[102]}
   );
   gpc1_1 gpc1_1_1521(
      {stage52[66]},
      {stage52[99]}
   );
   gpc1_1 gpc1_1_1522(
      {stage52[67]},
      {stage52[100]}
   );
   gpc1_1 gpc1_1_1523(
      {stage52[68]},
      {stage52[101]}
   );
   gpc1_1 gpc1_1_1524(
      {stage52[69]},
      {stage52[102]}
   );
   gpc1_1 gpc1_1_1525(
      {stage52[70]},
      {stage52[103]}
   );
   gpc1_1 gpc1_1_1526(
      {stage52[71]},
      {stage52[104]}
   );
   gpc1_1 gpc1_1_1527(
      {stage52[72]},
      {stage52[105]}
   );
   gpc1_1 gpc1_1_1528(
      {stage52[73]},
      {stage52[106]}
   );
   gpc606_5 gpc606_5_1529(
      {stage52[74], stage52[75], stage52[76], stage52[77], stage52[78], stage52[79]},
      {stage54[64], stage54[65], stage54[66], stage54[67], stage54[68], stage54[69]},
      {stage56[105], stage55[96], stage54[100], stage53[98], stage52[107]}
   );
   gpc606_5 gpc606_5_1530(
      {stage52[80], stage52[81], stage52[82], stage52[83], stage52[84], stage52[85]},
      {stage54[70], stage54[71], stage54[72], stage54[73], stage54[74], stage54[75]},
      {stage56[106], stage55[97], stage54[101], stage53[99], stage52[108]}
   );
   gpc606_5 gpc606_5_1531(
      {stage52[86], stage52[87], stage52[88], stage52[89], stage52[90], stage52[91]},
      {stage54[76], stage54[77], stage54[78], stage54[79], stage54[80], stage54[81]},
      {stage56[107], stage55[98], stage54[102], stage53[100], stage52[109]}
   );
   gpc1_1 gpc1_1_1532(
      {stage53[76]},
      {stage53[101]}
   );
   gpc1_1 gpc1_1_1533(
      {stage53[77]},
      {stage53[102]}
   );
   gpc1_1 gpc1_1_1534(
      {stage53[78]},
      {stage53[103]}
   );
   gpc1_1 gpc1_1_1535(
      {stage53[79]},
      {stage53[104]}
   );
   gpc1_1 gpc1_1_1536(
      {stage53[80]},
      {stage53[105]}
   );
   gpc1_1 gpc1_1_1537(
      {stage53[81]},
      {stage53[106]}
   );
   gpc1_1 gpc1_1_1538(
      {stage53[82]},
      {stage53[107]}
   );
   gpc1_1 gpc1_1_1539(
      {stage53[83]},
      {stage53[108]}
   );
   gpc1_1 gpc1_1_1540(
      {stage53[84]},
      {stage53[109]}
   );
   gpc615_5 gpc615_5_1541(
      {stage53[85], stage53[86], stage53[87], stage53[88], stage53[89]},
      {stage54[82]},
      {stage55[64], stage55[65], stage55[66], stage55[67], stage55[68], stage55[69]},
      {stage57[92], stage56[108], stage55[99], stage54[103], stage53[110]}
   );
   gpc615_5 gpc615_5_1542(
      {stage53[90], stage53[91], stage53[92], stage53[93], stage53[94]},
      {stage54[83]},
      {stage55[70], stage55[71], stage55[72], stage55[73], stage55[74], stage55[75]},
      {stage57[93], stage56[109], stage55[100], stage54[104], stage53[111]}
   );
   gpc1_1 gpc1_1_1543(
      {stage54[84]},
      {stage54[105]}
   );
   gpc1_1 gpc1_1_1544(
      {stage54[85]},
      {stage54[106]}
   );
   gpc1_1 gpc1_1_1545(
      {stage54[86]},
      {stage54[107]}
   );
   gpc1_1 gpc1_1_1546(
      {stage54[87]},
      {stage54[108]}
   );
   gpc1_1 gpc1_1_1547(
      {stage54[88]},
      {stage54[109]}
   );
   gpc1_1 gpc1_1_1548(
      {stage54[89]},
      {stage54[110]}
   );
   gpc1_1 gpc1_1_1549(
      {stage54[90]},
      {stage54[111]}
   );
   gpc1_1 gpc1_1_1550(
      {stage54[91]},
      {stage54[112]}
   );
   gpc1_1 gpc1_1_1551(
      {stage54[92]},
      {stage54[113]}
   );
   gpc615_5 gpc615_5_1552(
      {stage54[93], stage54[94], stage54[95], stage54[96], stage54[97]},
      {stage55[76]},
      {stage56[64], stage56[65], stage56[66], stage56[67], stage56[68], stage56[69]},
      {stage58[99], stage57[94], stage56[110], stage55[101], stage54[114]}
   );
   gpc1_1 gpc1_1_1553(
      {stage55[77]},
      {stage55[102]}
   );
   gpc1_1 gpc1_1_1554(
      {stage55[78]},
      {stage55[103]}
   );
   gpc615_5 gpc615_5_1555(
      {stage55[79], stage55[80], stage55[81], stage55[82], stage55[83]},
      {stage56[70]},
      {stage57[64], stage57[65], stage57[66], stage57[67], stage57[68], stage57[69]},
      {stage59[99], stage58[100], stage57[95], stage56[111], stage55[104]}
   );
   gpc615_5 gpc615_5_1556(
      {stage55[84], stage55[85], stage55[86], stage55[87], stage55[88]},
      {stage56[71]},
      {stage57[70], stage57[71], stage57[72], stage57[73], stage57[74], stage57[75]},
      {stage59[100], stage58[101], stage57[96], stage56[112], stage55[105]}
   );
   gpc615_5 gpc615_5_1557(
      {stage55[89], stage55[90], stage55[91], stage55[92], stage55[93]},
      {stage56[72]},
      {stage57[76], stage57[77], stage57[78], stage57[79], stage57[80], stage57[81]},
      {stage59[101], stage58[102], stage57[97], stage56[113], stage55[106]}
   );
   gpc1_1 gpc1_1_1558(
      {stage56[73]},
      {stage56[114]}
   );
   gpc1_1 gpc1_1_1559(
      {stage56[74]},
      {stage56[115]}
   );
   gpc1_1 gpc1_1_1560(
      {stage56[75]},
      {stage56[116]}
   );
   gpc1_1 gpc1_1_1561(
      {stage56[76]},
      {stage56[117]}
   );
   gpc1_1 gpc1_1_1562(
      {stage56[77]},
      {stage56[118]}
   );
   gpc1_1 gpc1_1_1563(
      {stage56[78]},
      {stage56[119]}
   );
   gpc1_1 gpc1_1_1564(
      {stage56[79]},
      {stage56[120]}
   );
   gpc1_1 gpc1_1_1565(
      {stage56[80]},
      {stage56[121]}
   );
   gpc1_1 gpc1_1_1566(
      {stage56[81]},
      {stage56[122]}
   );
   gpc1_1 gpc1_1_1567(
      {stage56[82]},
      {stage56[123]}
   );
   gpc1_1 gpc1_1_1568(
      {stage56[83]},
      {stage56[124]}
   );
   gpc1_1 gpc1_1_1569(
      {stage56[84]},
      {stage56[125]}
   );
   gpc615_5 gpc615_5_1570(
      {stage56[85], stage56[86], stage56[87], stage56[88], stage56[89]},
      {stage57[82]},
      {stage58[64], stage58[65], stage58[66], stage58[67], stage58[68], stage58[69]},
      {stage60[98], stage59[102], stage58[103], stage57[98], stage56[126]}
   );
   gpc615_5 gpc615_5_1571(
      {stage56[90], stage56[91], stage56[92], stage56[93], stage56[94]},
      {stage57[83]},
      {stage58[70], stage58[71], stage58[72], stage58[73], stage58[74], stage58[75]},
      {stage60[99], stage59[103], stage58[104], stage57[99], stage56[127]}
   );
   gpc615_5 gpc615_5_1572(
      {stage56[95], stage56[96], stage56[97], stage56[98], stage56[99]},
      {stage57[84]},
      {stage58[76], stage58[77], stage58[78], stage58[79], stage58[80], stage58[81]},
      {stage60[100], stage59[104], stage58[105], stage57[100], stage56[128]}
   );
   gpc615_5 gpc615_5_1573(
      {stage56[100], stage56[101], stage56[102], stage56[103], stage56[104]},
      {stage57[85]},
      {stage58[82], stage58[83], stage58[84], stage58[85], stage58[86], stage58[87]},
      {stage60[101], stage59[105], stage58[106], stage57[101], stage56[129]}
   );
   gpc1_1 gpc1_1_1574(
      {stage57[86]},
      {stage57[102]}
   );
   gpc1_1 gpc1_1_1575(
      {stage57[87]},
      {stage57[103]}
   );
   gpc1_1 gpc1_1_1576(
      {stage57[88]},
      {stage57[104]}
   );
   gpc1_1 gpc1_1_1577(
      {stage57[89]},
      {stage57[105]}
   );
   gpc1_1 gpc1_1_1578(
      {stage57[90]},
      {stage57[106]}
   );
   gpc1_1 gpc1_1_1579(
      {stage57[91]},
      {stage57[107]}
   );
   gpc1_1 gpc1_1_1580(
      {stage58[88]},
      {stage58[107]}
   );
   gpc1_1 gpc1_1_1581(
      {stage58[89]},
      {stage58[108]}
   );
   gpc1_1 gpc1_1_1582(
      {stage58[90]},
      {stage58[109]}
   );
   gpc1_1 gpc1_1_1583(
      {stage58[91]},
      {stage58[110]}
   );
   gpc1_1 gpc1_1_1584(
      {stage58[92]},
      {stage58[111]}
   );
   gpc1_1 gpc1_1_1585(
      {stage58[93]},
      {stage58[112]}
   );
   gpc615_5 gpc615_5_1586(
      {stage58[94], stage58[95], stage58[96], stage58[97], stage58[98]},
      {stage59[64]},
      {stage60[64], stage60[65], stage60[66], stage60[67], stage60[68], stage60[69]},
      {stage62[93], stage61[104], stage60[102], stage59[106], stage58[113]}
   );
   gpc1_1 gpc1_1_1587(
      {stage59[65]},
      {stage59[107]}
   );
   gpc1_1 gpc1_1_1588(
      {stage59[66]},
      {stage59[108]}
   );
   gpc1_1 gpc1_1_1589(
      {stage59[67]},
      {stage59[109]}
   );
   gpc1_1 gpc1_1_1590(
      {stage59[68]},
      {stage59[110]}
   );
   gpc1_1 gpc1_1_1591(
      {stage59[69]},
      {stage59[111]}
   );
   gpc1_1 gpc1_1_1592(
      {stage59[70]},
      {stage59[112]}
   );
   gpc1_1 gpc1_1_1593(
      {stage59[71]},
      {stage59[113]}
   );
   gpc1_1 gpc1_1_1594(
      {stage59[72]},
      {stage59[114]}
   );
   gpc1_1 gpc1_1_1595(
      {stage59[73]},
      {stage59[115]}
   );
   gpc2135_5 gpc2135_5_1596(
      {stage59[74], stage59[75], stage59[76], stage59[77], stage59[78]},
      {stage60[70], stage60[71], stage60[72]},
      {stage61[64]},
      {stage62[64], stage62[65]},
      {stage63[97], stage62[94], stage61[105], stage60[103], stage59[116]}
   );
   gpc2135_5 gpc2135_5_1597(
      {stage59[79], stage59[80], stage59[81], stage59[82], stage59[83]},
      {stage60[73], stage60[74], stage60[75]},
      {stage61[65]},
      {stage62[66], stage62[67]},
      {stage63[98], stage62[95], stage61[106], stage60[104], stage59[117]}
   );
   gpc2135_5 gpc2135_5_1598(
      {stage59[84], stage59[85], stage59[86], stage59[87], stage59[88]},
      {stage60[76], stage60[77], stage60[78]},
      {stage61[66]},
      {stage62[68], stage62[69]},
      {stage63[99], stage62[96], stage61[107], stage60[105], stage59[118]}
   );
   gpc2135_5 gpc2135_5_1599(
      {stage59[89], stage59[90], stage59[91], stage59[92], stage59[93]},
      {stage60[79], stage60[80], stage60[81]},
      {stage61[67]},
      {stage62[70], stage62[71]},
      {stage63[100], stage62[97], stage61[108], stage60[106], stage59[119]}
   );
   gpc2135_5 gpc2135_5_1600(
      {stage59[94], stage59[95], stage59[96], stage59[97], stage59[98]},
      {stage60[82], stage60[83], stage60[84]},
      {stage61[68]},
      {stage62[72], stage62[73]},
      {stage63[101], stage62[98], stage61[109], stage60[107], stage59[120]}
   );
   gpc1_1 gpc1_1_1601(
      {stage60[85]},
      {stage60[108]}
   );
   gpc1_1 gpc1_1_1602(
      {stage60[86]},
      {stage60[109]}
   );
   gpc1_1 gpc1_1_1603(
      {stage60[87]},
      {stage60[110]}
   );
   gpc1_1 gpc1_1_1604(
      {stage60[88]},
      {stage60[111]}
   );
   gpc1_1 gpc1_1_1605(
      {stage60[89]},
      {stage60[112]}
   );
   gpc1_1 gpc1_1_1606(
      {stage60[90]},
      {stage60[113]}
   );
   gpc1_1 gpc1_1_1607(
      {stage60[91]},
      {stage60[114]}
   );
   gpc1_1 gpc1_1_1608(
      {stage60[92]},
      {stage60[115]}
   );
   gpc615_5 gpc615_5_1609(
      {stage60[93], stage60[94], stage60[95], stage60[96], stage60[97]},
      {stage61[69]},
      {stage62[74], stage62[75], stage62[76], stage62[77], stage62[78], stage62[79]},
      {stage64[16], stage63[102], stage62[99], stage61[110], stage60[116]}
   );
   gpc1_1 gpc1_1_1610(
      {stage61[70]},
      {stage61[111]}
   );
   gpc1_1 gpc1_1_1611(
      {stage61[71]},
      {stage61[112]}
   );
   gpc1_1 gpc1_1_1612(
      {stage61[72]},
      {stage61[113]}
   );
   gpc1_1 gpc1_1_1613(
      {stage61[73]},
      {stage61[114]}
   );
   gpc1_1 gpc1_1_1614(
      {stage61[74]},
      {stage61[115]}
   );
   gpc1_1 gpc1_1_1615(
      {stage61[75]},
      {stage61[116]}
   );
   gpc1_1 gpc1_1_1616(
      {stage61[76]},
      {stage61[117]}
   );
   gpc1_1 gpc1_1_1617(
      {stage61[77]},
      {stage61[118]}
   );
   gpc1_1 gpc1_1_1618(
      {stage61[78]},
      {stage61[119]}
   );
   gpc1_1 gpc1_1_1619(
      {stage61[79]},
      {stage61[120]}
   );
   gpc606_5 gpc606_5_1620(
      {stage61[80], stage61[81], stage61[82], stage61[83], stage61[84], stage61[85]},
      {stage63[64], stage63[65], stage63[66], stage63[67], stage63[68], stage63[69]},
      {stage65[8], stage64[17], stage63[103], stage62[100], stage61[121]}
   );
   gpc606_5 gpc606_5_1621(
      {stage61[86], stage61[87], stage61[88], stage61[89], stage61[90], stage61[91]},
      {stage63[70], stage63[71], stage63[72], stage63[73], stage63[74], stage63[75]},
      {stage65[9], stage64[18], stage63[104], stage62[101], stage61[122]}
   );
   gpc606_5 gpc606_5_1622(
      {stage61[92], stage61[93], stage61[94], stage61[95], stage61[96], stage61[97]},
      {stage63[76], stage63[77], stage63[78], stage63[79], stage63[80], stage63[81]},
      {stage65[10], stage64[19], stage63[105], stage62[102], stage61[123]}
   );
   gpc606_5 gpc606_5_1623(
      {stage61[98], stage61[99], stage61[100], stage61[101], stage61[102], stage61[103]},
      {stage63[82], stage63[83], stage63[84], stage63[85], stage63[86], stage63[87]},
      {stage65[11], stage64[20], stage63[106], stage62[103], stage61[124]}
   );
   gpc1_1 gpc1_1_1624(
      {stage62[80]},
      {stage62[104]}
   );
   gpc1_1 gpc1_1_1625(
      {stage62[81]},
      {stage62[105]}
   );
   gpc1_1 gpc1_1_1626(
      {stage62[82]},
      {stage62[106]}
   );
   gpc1_1 gpc1_1_1627(
      {stage62[83]},
      {stage62[107]}
   );
   gpc606_5 gpc606_5_1628(
      {stage62[84], stage62[85], stage62[86], stage62[87], stage62[88], stage62[89]},
      {stage64[0], stage64[1], stage64[2], stage64[3], stage64[4], stage64[5]},
      {stage66[0], stage65[12], stage64[21], stage63[107], stage62[108]}
   );
   gpc1343_5 gpc1343_5_1629(
      {stage62[90], stage62[91], stage62[92]},
      {stage63[88], stage63[89], stage63[90], stage63[91]},
      {stage64[6], stage64[7], stage64[8]},
      {stage65[0]},
      {stage66[1], stage65[13], stage64[22], stage63[108], stage62[109]}
   );
   gpc606_5 gpc606_5_1630(
      {stage63[92], stage63[93], stage63[94], stage63[95], stage63[96], 1'h0},
      {stage65[1], stage65[2], stage65[3], stage65[4], stage65[5], stage65[6]},
      {stage67[0], stage66[2], stage65[14], stage64[23], stage63[109]}
   );
   gpc1_1 gpc1_1_1631(
      {stage64[9]},
      {stage64[24]}
   );
   gpc1_1 gpc1_1_1632(
      {stage64[10]},
      {stage64[25]}
   );
   gpc1_1 gpc1_1_1633(
      {stage64[11]},
      {stage64[26]}
   );
   gpc1_1 gpc1_1_1634(
      {stage64[12]},
      {stage64[27]}
   );
   gpc1_1 gpc1_1_1635(
      {stage64[13]},
      {stage64[28]}
   );
   gpc1_1 gpc1_1_1636(
      {stage64[14]},
      {stage64[29]}
   );
   gpc1_1 gpc1_1_1637(
      {stage64[15]},
      {stage64[30]}
   );
   gpc1_1 gpc1_1_1638(
      {stage65[7]},
      {stage65[15]}
   );
   gpc1_1 gpc1_1_1639(
      {stage00[80]},
      {stage00[86]}
   );
   gpc1_1 gpc1_1_1640(
      {stage00[81]},
      {stage00[87]}
   );
   gpc1_1 gpc1_1_1641(
      {stage00[82]},
      {stage00[88]}
   );
   gpc1_1 gpc1_1_1642(
      {stage00[83]},
      {stage00[89]}
   );
   gpc1_1 gpc1_1_1643(
      {stage00[84]},
      {stage00[90]}
   );
   gpc1_1 gpc1_1_1644(
      {stage00[85]},
      {stage00[91]}
   );
   gpc1_1 gpc1_1_1645(
      {stage01[110]},
      {stage01[123]}
   );
   gpc606_5 gpc606_5_1646(
      {stage01[111], stage01[112], stage01[113], stage01[114], stage01[115], stage01[116]},
      {stage03[121], stage03[122], stage03[123], stage03[124], stage03[125], stage03[126]},
      {stage05[111], stage04[112], stage03[133], stage02[105], stage01[124]}
   );
   gpc606_5 gpc606_5_1647(
      {stage01[117], stage01[118], stage01[119], stage01[120], stage01[121], stage01[122]},
      {stage03[127], stage03[128], stage03[129], stage03[130], stage03[131], stage03[132]},
      {stage05[112], stage04[113], stage03[134], stage02[106], stage01[125]}
   );
   gpc1_1 gpc1_1_1648(
      {stage02[86]},
      {stage02[107]}
   );
   gpc606_5 gpc606_5_1649(
      {stage02[87], stage02[88], stage02[89], stage02[90], stage02[91], stage02[92]},
      {stage04[93], stage04[94], stage04[95], stage04[96], stage04[97], stage04[98]},
      {stage06[99], stage05[113], stage04[114], stage03[135], stage02[108]}
   );
   gpc606_5 gpc606_5_1650(
      {stage02[93], stage02[94], stage02[95], stage02[96], stage02[97], stage02[98]},
      {stage04[99], stage04[100], stage04[101], stage04[102], stage04[103], stage04[104]},
      {stage06[100], stage05[114], stage04[115], stage03[136], stage02[109]}
   );
   gpc606_5 gpc606_5_1651(
      {stage02[99], stage02[100], stage02[101], stage02[102], stage02[103], stage02[104]},
      {stage04[105], stage04[106], stage04[107], stage04[108], stage04[109], stage04[110]},
      {stage06[101], stage05[115], stage04[116], stage03[137], stage02[110]}
   );
   gpc1_1 gpc1_1_1652(
      {stage04[111]},
      {stage04[117]}
   );
   gpc1_1 gpc1_1_1653(
      {stage05[90]},
      {stage05[116]}
   );
   gpc1_1 gpc1_1_1654(
      {stage05[91]},
      {stage05[117]}
   );
   gpc1_1 gpc1_1_1655(
      {stage05[92]},
      {stage05[118]}
   );
   gpc606_5 gpc606_5_1656(
      {stage05[93], stage05[94], stage05[95], stage05[96], stage05[97], stage05[98]},
      {stage07[97], stage07[98], stage07[99], stage07[100], stage07[101], stage07[102]},
      {stage09[152], stage08[119], stage07[111], stage06[102], stage05[119]}
   );
   gpc606_5 gpc606_5_1657(
      {stage05[99], stage05[100], stage05[101], stage05[102], stage05[103], stage05[104]},
      {stage07[103], stage07[104], stage07[105], stage07[106], stage07[107], stage07[108]},
      {stage09[153], stage08[120], stage07[112], stage06[103], stage05[120]}
   );
   gpc606_5 gpc606_5_1658(
      {stage05[105], stage05[106], stage05[107], stage05[108], stage05[109], stage05[110]},
      {stage07[109], stage07[110], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage09[154], stage08[121], stage07[113], stage06[104], stage05[121]}
   );
   gpc1_1 gpc1_1_1659(
      {stage06[90]},
      {stage06[105]}
   );
   gpc1_1 gpc1_1_1660(
      {stage06[91]},
      {stage06[106]}
   );
   gpc1_1 gpc1_1_1661(
      {stage06[92]},
      {stage06[107]}
   );
   gpc606_5 gpc606_5_1662(
      {stage06[93], stage06[94], stage06[95], stage06[96], stage06[97], stage06[98]},
      {stage08[102], stage08[103], stage08[104], stage08[105], stage08[106], stage08[107]},
      {stage10[130], stage09[155], stage08[122], stage07[114], stage06[108]}
   );
   gpc606_5 gpc606_5_1663(
      {stage08[108], stage08[109], stage08[110], stage08[111], stage08[112], stage08[113]},
      {stage10[110], stage10[111], stage10[112], stage10[113], stage10[114], stage10[115]},
      {stage12[131], stage11[134], stage10[131], stage09[156], stage08[123]}
   );
   gpc606_5 gpc606_5_1664(
      {stage08[114], stage08[115], stage08[116], stage08[117], stage08[118], 1'h0},
      {stage10[116], stage10[117], stage10[118], stage10[119], stage10[120], stage10[121]},
      {stage12[132], stage11[135], stage10[132], stage09[157], stage08[124]}
   );
   gpc1_1 gpc1_1_1665(
      {stage09[123]},
      {stage09[158]}
   );
   gpc1_1 gpc1_1_1666(
      {stage09[124]},
      {stage09[159]}
   );
   gpc1_1 gpc1_1_1667(
      {stage09[125]},
      {stage09[160]}
   );
   gpc1_1 gpc1_1_1668(
      {stage09[126]},
      {stage09[161]}
   );
   gpc1_1 gpc1_1_1669(
      {stage09[127]},
      {stage09[162]}
   );
   gpc606_5 gpc606_5_1670(
      {stage09[128], stage09[129], stage09[130], stage09[131], stage09[132], stage09[133]},
      {stage11[93], stage11[94], stage11[95], stage11[96], stage11[97], stage11[98]},
      {stage13[107], stage12[133], stage11[136], stage10[133], stage09[163]}
   );
   gpc606_5 gpc606_5_1671(
      {stage09[134], stage09[135], stage09[136], stage09[137], stage09[138], stage09[139]},
      {stage11[99], stage11[100], stage11[101], stage11[102], stage11[103], stage11[104]},
      {stage13[108], stage12[134], stage11[137], stage10[134], stage09[164]}
   );
   gpc606_5 gpc606_5_1672(
      {stage09[140], stage09[141], stage09[142], stage09[143], stage09[144], stage09[145]},
      {stage11[105], stage11[106], stage11[107], stage11[108], stage11[109], stage11[110]},
      {stage13[109], stage12[135], stage11[138], stage10[135], stage09[165]}
   );
   gpc606_5 gpc606_5_1673(
      {stage09[146], stage09[147], stage09[148], stage09[149], stage09[150], stage09[151]},
      {stage11[111], stage11[112], stage11[113], stage11[114], stage11[115], stage11[116]},
      {stage13[110], stage12[136], stage11[139], stage10[136], stage09[166]}
   );
   gpc615_5 gpc615_5_1674(
      {stage10[122], stage10[123], stage10[124], stage10[125], stage10[126]},
      {stage11[117]},
      {stage12[110], stage12[111], stage12[112], stage12[113], stage12[114], stage12[115]},
      {stage14[105], stage13[111], stage12[137], stage11[140], stage10[137]}
   );
   gpc615_5 gpc615_5_1675(
      {stage10[127], stage10[128], stage10[129], 1'h0, 1'h0},
      {stage11[118]},
      {stage12[116], stage12[117], stage12[118], stage12[119], stage12[120], stage12[121]},
      {stage14[106], stage13[112], stage12[138], stage11[141], stage10[138]}
   );
   gpc1_1 gpc1_1_1676(
      {stage11[119]},
      {stage11[142]}
   );
   gpc1_1 gpc1_1_1677(
      {stage11[120]},
      {stage11[143]}
   );
   gpc1_1 gpc1_1_1678(
      {stage11[121]},
      {stage11[144]}
   );
   gpc1_1 gpc1_1_1679(
      {stage11[122]},
      {stage11[145]}
   );
   gpc1_1 gpc1_1_1680(
      {stage11[123]},
      {stage11[146]}
   );
   gpc1_1 gpc1_1_1681(
      {stage11[124]},
      {stage11[147]}
   );
   gpc1_1 gpc1_1_1682(
      {stage11[125]},
      {stage11[148]}
   );
   gpc1_1 gpc1_1_1683(
      {stage11[126]},
      {stage11[149]}
   );
   gpc1_1 gpc1_1_1684(
      {stage11[127]},
      {stage11[150]}
   );
   gpc1_1 gpc1_1_1685(
      {stage11[128]},
      {stage11[151]}
   );
   gpc615_5 gpc615_5_1686(
      {stage11[129], stage11[130], stage11[131], stage11[132], stage11[133]},
      {stage12[122]},
      {stage13[90], stage13[91], stage13[92], stage13[93], stage13[94], stage13[95]},
      {stage15[145], stage14[107], stage13[113], stage12[139], stage11[152]}
   );
   gpc1_1 gpc1_1_1687(
      {stage12[123]},
      {stage12[140]}
   );
   gpc1_1 gpc1_1_1688(
      {stage12[124]},
      {stage12[141]}
   );
   gpc606_5 gpc606_5_1689(
      {stage12[125], stage12[126], stage12[127], stage12[128], stage12[129], stage12[130]},
      {stage14[94], stage14[95], stage14[96], stage14[97], stage14[98], stage14[99]},
      {stage16[105], stage15[146], stage14[108], stage13[114], stage12[142]}
   );
   gpc1_1 gpc1_1_1690(
      {stage13[96]},
      {stage13[115]}
   );
   gpc1_1 gpc1_1_1691(
      {stage13[97]},
      {stage13[116]}
   );
   gpc1_1 gpc1_1_1692(
      {stage13[98]},
      {stage13[117]}
   );
   gpc1_1 gpc1_1_1693(
      {stage13[99]},
      {stage13[118]}
   );
   gpc1_1 gpc1_1_1694(
      {stage13[100]},
      {stage13[119]}
   );
   gpc1_1 gpc1_1_1695(
      {stage13[101]},
      {stage13[120]}
   );
   gpc1_1 gpc1_1_1696(
      {stage13[102]},
      {stage13[121]}
   );
   gpc1_1 gpc1_1_1697(
      {stage13[103]},
      {stage13[122]}
   );
   gpc1_1 gpc1_1_1698(
      {stage13[104]},
      {stage13[123]}
   );
   gpc1_1 gpc1_1_1699(
      {stage13[105]},
      {stage13[124]}
   );
   gpc1_1 gpc1_1_1700(
      {stage13[106]},
      {stage13[125]}
   );
   gpc615_5 gpc615_5_1701(
      {stage14[100], stage14[101], stage14[102], stage14[103], stage14[104]},
      {stage15[124]},
      {stage16[90], stage16[91], stage16[92], stage16[93], stage16[94], stage16[95]},
      {stage18[102], stage17[138], stage16[106], stage15[147], stage14[109]}
   );
   gpc1_1 gpc1_1_1702(
      {stage15[125]},
      {stage15[148]}
   );
   gpc1_1 gpc1_1_1703(
      {stage15[126]},
      {stage15[149]}
   );
   gpc1_1 gpc1_1_1704(
      {stage15[127]},
      {stage15[150]}
   );
   gpc1_1 gpc1_1_1705(
      {stage15[128]},
      {stage15[151]}
   );
   gpc1_1 gpc1_1_1706(
      {stage15[129]},
      {stage15[152]}
   );
   gpc615_5 gpc615_5_1707(
      {stage15[130], stage15[131], stage15[132], stage15[133], stage15[134]},
      {stage16[96]},
      {stage17[104], stage17[105], stage17[106], stage17[107], stage17[108], stage17[109]},
      {stage19[115], stage18[103], stage17[139], stage16[107], stage15[153]}
   );
   gpc615_5 gpc615_5_1708(
      {stage15[135], stage15[136], stage15[137], stage15[138], stage15[139]},
      {stage16[97]},
      {stage17[110], stage17[111], stage17[112], stage17[113], stage17[114], stage17[115]},
      {stage19[116], stage18[104], stage17[140], stage16[108], stage15[154]}
   );
   gpc615_5 gpc615_5_1709(
      {stage15[140], stage15[141], stage15[142], stage15[143], stage15[144]},
      {stage16[98]},
      {stage17[116], stage17[117], stage17[118], stage17[119], stage17[120], stage17[121]},
      {stage19[117], stage18[105], stage17[141], stage16[109], stage15[155]}
   );
   gpc606_5 gpc606_5_1710(
      {stage16[99], stage16[100], stage16[101], stage16[102], stage16[103], stage16[104]},
      {stage18[85], stage18[86], stage18[87], stage18[88], stage18[89], stage18[90]},
      {stage20[125], stage19[118], stage18[106], stage17[142], stage16[110]}
   );
   gpc1_1 gpc1_1_1711(
      {stage17[122]},
      {stage17[143]}
   );
   gpc1_1 gpc1_1_1712(
      {stage17[123]},
      {stage17[144]}
   );
   gpc1_1 gpc1_1_1713(
      {stage17[124]},
      {stage17[145]}
   );
   gpc1_1 gpc1_1_1714(
      {stage17[125]},
      {stage17[146]}
   );
   gpc606_5 gpc606_5_1715(
      {stage17[126], stage17[127], stage17[128], stage17[129], stage17[130], stage17[131]},
      {stage19[99], stage19[100], stage19[101], stage19[102], stage19[103], stage19[104]},
      {stage21[105], stage20[126], stage19[119], stage18[107], stage17[147]}
   );
   gpc606_5 gpc606_5_1716(
      {stage17[132], stage17[133], stage17[134], stage17[135], stage17[136], stage17[137]},
      {stage19[105], stage19[106], stage19[107], stage19[108], stage19[109], stage19[110]},
      {stage21[106], stage20[127], stage19[120], stage18[108], stage17[148]}
   );
   gpc1_1 gpc1_1_1717(
      {stage18[91]},
      {stage18[109]}
   );
   gpc1_1 gpc1_1_1718(
      {stage18[92]},
      {stage18[110]}
   );
   gpc1_1 gpc1_1_1719(
      {stage18[93]},
      {stage18[111]}
   );
   gpc1_1 gpc1_1_1720(
      {stage18[94]},
      {stage18[112]}
   );
   gpc1_1 gpc1_1_1721(
      {stage18[95]},
      {stage18[113]}
   );
   gpc1_1 gpc1_1_1722(
      {stage18[96]},
      {stage18[114]}
   );
   gpc1_1 gpc1_1_1723(
      {stage18[97]},
      {stage18[115]}
   );
   gpc1_1 gpc1_1_1724(
      {stage18[98]},
      {stage18[116]}
   );
   gpc1_1 gpc1_1_1725(
      {stage18[99]},
      {stage18[117]}
   );
   gpc1_1 gpc1_1_1726(
      {stage18[100]},
      {stage18[118]}
   );
   gpc1_1 gpc1_1_1727(
      {stage18[101]},
      {stage18[119]}
   );
   gpc615_5 gpc615_5_1728(
      {stage19[111], stage19[112], stage19[113], stage19[114], 1'h0},
      {stage20[106]},
      {stage21[91], stage21[92], stage21[93], stage21[94], stage21[95], stage21[96]},
      {stage23[119], stage22[109], stage21[107], stage20[128], stage19[121]}
   );
   gpc1_1 gpc1_1_1729(
      {stage20[107]},
      {stage20[129]}
   );
   gpc1_1 gpc1_1_1730(
      {stage20[108]},
      {stage20[130]}
   );
   gpc1_1 gpc1_1_1731(
      {stage20[109]},
      {stage20[131]}
   );
   gpc1_1 gpc1_1_1732(
      {stage20[110]},
      {stage20[132]}
   );
   gpc1_1 gpc1_1_1733(
      {stage20[111]},
      {stage20[133]}
   );
   gpc1_1 gpc1_1_1734(
      {stage20[112]},
      {stage20[134]}
   );
   gpc1_1 gpc1_1_1735(
      {stage20[113]},
      {stage20[135]}
   );
   gpc1_1 gpc1_1_1736(
      {stage20[114]},
      {stage20[136]}
   );
   gpc1_1 gpc1_1_1737(
      {stage20[115]},
      {stage20[137]}
   );
   gpc1_1 gpc1_1_1738(
      {stage20[116]},
      {stage20[138]}
   );
   gpc1_1 gpc1_1_1739(
      {stage20[117]},
      {stage20[139]}
   );
   gpc1_1 gpc1_1_1740(
      {stage20[118]},
      {stage20[140]}
   );
   gpc1_1 gpc1_1_1741(
      {stage20[119]},
      {stage20[141]}
   );
   gpc1_1 gpc1_1_1742(
      {stage20[120]},
      {stage20[142]}
   );
   gpc1_1 gpc1_1_1743(
      {stage20[121]},
      {stage20[143]}
   );
   gpc1_1 gpc1_1_1744(
      {stage20[122]},
      {stage20[144]}
   );
   gpc1_1 gpc1_1_1745(
      {stage20[123]},
      {stage20[145]}
   );
   gpc1_1 gpc1_1_1746(
      {stage20[124]},
      {stage20[146]}
   );
   gpc1_1 gpc1_1_1747(
      {stage21[97]},
      {stage21[108]}
   );
   gpc1_1 gpc1_1_1748(
      {stage21[98]},
      {stage21[109]}
   );
   gpc1_1 gpc1_1_1749(
      {stage21[99]},
      {stage21[110]}
   );
   gpc615_5 gpc615_5_1750(
      {stage21[100], stage21[101], stage21[102], stage21[103], stage21[104]},
      {stage22[99]},
      {stage23[95], stage23[96], stage23[97], stage23[98], stage23[99], stage23[100]},
      {stage25[117], stage24[112], stage23[120], stage22[110], stage21[111]}
   );
   gpc1415_5 gpc1415_5_1751(
      {stage22[100], stage22[101], stage22[102], stage22[103], stage22[104]},
      {stage23[101]},
      {stage24[98], stage24[99], stage24[100], stage24[101]},
      {stage25[98]},
      {stage26[96], stage25[118], stage24[113], stage23[121], stage22[111]}
   );
   gpc1415_5 gpc1415_5_1752(
      {stage22[105], stage22[106], stage22[107], stage22[108], 1'h0},
      {stage23[102]},
      {stage24[102], stage24[103], stage24[104], stage24[105]},
      {stage25[99]},
      {stage26[97], stage25[119], stage24[114], stage23[122], stage22[112]}
   );
   gpc1_1 gpc1_1_1753(
      {stage23[103]},
      {stage23[123]}
   );
   gpc1_1 gpc1_1_1754(
      {stage23[104]},
      {stage23[124]}
   );
   gpc1_1 gpc1_1_1755(
      {stage23[105]},
      {stage23[125]}
   );
   gpc1_1 gpc1_1_1756(
      {stage23[106]},
      {stage23[126]}
   );
   gpc1_1 gpc1_1_1757(
      {stage23[107]},
      {stage23[127]}
   );
   gpc1_1 gpc1_1_1758(
      {stage23[108]},
      {stage23[128]}
   );
   gpc1_1 gpc1_1_1759(
      {stage23[109]},
      {stage23[129]}
   );
   gpc1_1 gpc1_1_1760(
      {stage23[110]},
      {stage23[130]}
   );
   gpc1_1 gpc1_1_1761(
      {stage23[111]},
      {stage23[131]}
   );
   gpc1_1 gpc1_1_1762(
      {stage23[112]},
      {stage23[132]}
   );
   gpc1_1 gpc1_1_1763(
      {stage23[113]},
      {stage23[133]}
   );
   gpc615_5 gpc615_5_1764(
      {stage23[114], stage23[115], stage23[116], stage23[117], stage23[118]},
      {stage24[106]},
      {stage25[100], stage25[101], stage25[102], stage25[103], stage25[104], stage25[105]},
      {stage27[127], stage26[98], stage25[120], stage24[115], stage23[134]}
   );
   gpc615_5 gpc615_5_1765(
      {stage24[107], stage24[108], stage24[109], stage24[110], stage24[111]},
      {stage25[106]},
      {stage26[87], stage26[88], stage26[89], stage26[90], stage26[91], stage26[92]},
      {stage28[125], stage27[128], stage26[99], stage25[121], stage24[116]}
   );
   gpc1_1 gpc1_1_1766(
      {stage25[107]},
      {stage25[122]}
   );
   gpc1_1 gpc1_1_1767(
      {stage25[108]},
      {stage25[123]}
   );
   gpc1_1 gpc1_1_1768(
      {stage25[109]},
      {stage25[124]}
   );
   gpc1_1 gpc1_1_1769(
      {stage25[110]},
      {stage25[125]}
   );
   gpc1_1 gpc1_1_1770(
      {stage25[111]},
      {stage25[126]}
   );
   gpc1_1 gpc1_1_1771(
      {stage25[112]},
      {stage25[127]}
   );
   gpc1_1 gpc1_1_1772(
      {stage25[113]},
      {stage25[128]}
   );
   gpc1_1 gpc1_1_1773(
      {stage25[114]},
      {stage25[129]}
   );
   gpc1_1 gpc1_1_1774(
      {stage25[115]},
      {stage25[130]}
   );
   gpc1_1 gpc1_1_1775(
      {stage25[116]},
      {stage25[131]}
   );
   gpc1_1 gpc1_1_1776(
      {stage26[93]},
      {stage26[100]}
   );
   gpc1_1 gpc1_1_1777(
      {stage26[94]},
      {stage26[101]}
   );
   gpc1_1 gpc1_1_1778(
      {stage26[95]},
      {stage26[102]}
   );
   gpc1_1 gpc1_1_1779(
      {stage27[104]},
      {stage27[129]}
   );
   gpc1_1 gpc1_1_1780(
      {stage27[105]},
      {stage27[130]}
   );
   gpc1_1 gpc1_1_1781(
      {stage27[106]},
      {stage27[131]}
   );
   gpc2135_5 gpc2135_5_1782(
      {stage27[107], stage27[108], stage27[109], stage27[110], stage27[111]},
      {stage28[90], stage28[91], stage28[92]},
      {stage29[94]},
      {stage30[94], stage30[95]},
      {stage31[107], stage30[121], stage29[99], stage28[126], stage27[132]}
   );
   gpc2135_5 gpc2135_5_1783(
      {stage27[112], stage27[113], stage27[114], stage27[115], stage27[116]},
      {stage28[93], stage28[94], stage28[95]},
      {stage29[95]},
      {stage30[96], stage30[97]},
      {stage31[108], stage30[122], stage29[100], stage28[127], stage27[133]}
   );
   gpc2135_5 gpc2135_5_1784(
      {stage27[117], stage27[118], stage27[119], stage27[120], stage27[121]},
      {stage28[96], stage28[97], stage28[98]},
      {stage29[96]},
      {stage30[98], stage30[99]},
      {stage31[109], stage30[123], stage29[101], stage28[128], stage27[134]}
   );
   gpc2135_5 gpc2135_5_1785(
      {stage27[122], stage27[123], stage27[124], stage27[125], stage27[126]},
      {stage28[99], stage28[100], stage28[101]},
      {stage29[97]},
      {stage30[100], stage30[101]},
      {stage31[110], stage30[124], stage29[102], stage28[129], stage27[135]}
   );
   gpc1_1 gpc1_1_1786(
      {stage28[102]},
      {stage28[130]}
   );
   gpc1_1 gpc1_1_1787(
      {stage28[103]},
      {stage28[131]}
   );
   gpc1_1 gpc1_1_1788(
      {stage28[104]},
      {stage28[132]}
   );
   gpc1_1 gpc1_1_1789(
      {stage28[105]},
      {stage28[133]}
   );
   gpc1_1 gpc1_1_1790(
      {stage28[106]},
      {stage28[134]}
   );
   gpc606_5 gpc606_5_1791(
      {stage28[107], stage28[108], stage28[109], stage28[110], stage28[111], stage28[112]},
      {stage30[102], stage30[103], stage30[104], stage30[105], stage30[106], stage30[107]},
      {stage32[105], stage31[111], stage30[125], stage29[103], stage28[135]}
   );
   gpc606_5 gpc606_5_1792(
      {stage28[113], stage28[114], stage28[115], stage28[116], stage28[117], stage28[118]},
      {stage30[108], stage30[109], stage30[110], stage30[111], stage30[112], stage30[113]},
      {stage32[106], stage31[112], stage30[126], stage29[104], stage28[136]}
   );
   gpc606_5 gpc606_5_1793(
      {stage28[119], stage28[120], stage28[121], stage28[122], stage28[123], stage28[124]},
      {stage30[114], stage30[115], stage30[116], stage30[117], stage30[118], stage30[119]},
      {stage32[107], stage31[113], stage30[127], stage29[105], stage28[137]}
   );
   gpc1_1 gpc1_1_1794(
      {stage29[98]},
      {stage29[106]}
   );
   gpc615_5 gpc615_5_1795(
      {stage30[120], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage31[91]},
      {stage32[97], stage32[98], stage32[99], stage32[100], stage32[101], stage32[102]},
      {stage34[102], stage33[106], stage32[108], stage31[114], stage30[128]}
   );
   gpc1_1 gpc1_1_1796(
      {stage31[92]},
      {stage31[115]}
   );
   gpc1_1 gpc1_1_1797(
      {stage31[93]},
      {stage31[116]}
   );
   gpc1_1 gpc1_1_1798(
      {stage31[94]},
      {stage31[117]}
   );
   gpc1_1 gpc1_1_1799(
      {stage31[95]},
      {stage31[118]}
   );
   gpc1_1 gpc1_1_1800(
      {stage31[96]},
      {stage31[119]}
   );
   gpc615_5 gpc615_5_1801(
      {stage31[97], stage31[98], stage31[99], stage31[100], stage31[101]},
      {stage32[103]},
      {stage33[90], stage33[91], stage33[92], stage33[93], stage33[94], stage33[95]},
      {stage35[106], stage34[103], stage33[107], stage32[109], stage31[120]}
   );
   gpc615_5 gpc615_5_1802(
      {stage31[102], stage31[103], stage31[104], stage31[105], stage31[106]},
      {stage32[104]},
      {stage33[96], stage33[97], stage33[98], stage33[99], stage33[100], stage33[101]},
      {stage35[107], stage34[104], stage33[108], stage32[110], stage31[121]}
   );
   gpc606_5 gpc606_5_1803(
      {stage33[102], stage33[103], stage33[104], stage33[105], 1'h0, 1'h0},
      {stage35[91], stage35[92], stage35[93], stage35[94], stage35[95], stage35[96]},
      {stage37[109], stage36[121], stage35[108], stage34[105], stage33[109]}
   );
   gpc135_4 gpc135_4_1804(
      {stage34[88], stage34[89], stage34[90], stage34[91], stage34[92]},
      {stage35[97], stage35[98], stage35[99]},
      {stage36[107]},
      {stage37[110], stage36[122], stage35[109], stage34[106]}
   );
   gpc135_4 gpc135_4_1805(
      {stage34[93], stage34[94], stage34[95], stage34[96], stage34[97]},
      {stage35[100], stage35[101], stage35[102]},
      {stage36[108]},
      {stage37[111], stage36[123], stage35[110], stage34[107]}
   );
   gpc135_4 gpc135_4_1806(
      {stage34[98], stage34[99], stage34[100], stage34[101], 1'h0},
      {stage35[103], stage35[104], stage35[105]},
      {stage36[109]},
      {stage37[112], stage36[124], stage35[111], stage34[108]}
   );
   gpc1_1 gpc1_1_1807(
      {stage36[110]},
      {stage36[125]}
   );
   gpc1_1 gpc1_1_1808(
      {stage36[111]},
      {stage36[126]}
   );
   gpc1_1 gpc1_1_1809(
      {stage36[112]},
      {stage36[127]}
   );
   gpc1_1 gpc1_1_1810(
      {stage36[113]},
      {stage36[128]}
   );
   gpc1_1 gpc1_1_1811(
      {stage36[114]},
      {stage36[129]}
   );
   gpc1343_5 gpc1343_5_1812(
      {stage36[115], stage36[116], stage36[117]},
      {stage37[96], stage37[97], stage37[98], stage37[99]},
      {stage38[88], stage38[89], stage38[90]},
      {stage39[92]},
      {stage40[120], stage39[104], stage38[105], stage37[113], stage36[130]}
   );
   gpc1343_5 gpc1343_5_1813(
      {stage36[118], stage36[119], stage36[120]},
      {stage37[100], stage37[101], stage37[102], stage37[103]},
      {stage38[91], stage38[92], stage38[93]},
      {stage39[93]},
      {stage40[121], stage39[105], stage38[106], stage37[114], stage36[131]}
   );
   gpc1_1 gpc1_1_1814(
      {stage37[104]},
      {stage37[115]}
   );
   gpc1_1 gpc1_1_1815(
      {stage37[105]},
      {stage37[116]}
   );
   gpc1_1 gpc1_1_1816(
      {stage37[106]},
      {stage37[117]}
   );
   gpc1_1 gpc1_1_1817(
      {stage37[107]},
      {stage37[118]}
   );
   gpc1_1 gpc1_1_1818(
      {stage37[108]},
      {stage37[119]}
   );
   gpc1_1 gpc1_1_1819(
      {stage38[94]},
      {stage38[107]}
   );
   gpc1_1 gpc1_1_1820(
      {stage38[95]},
      {stage38[108]}
   );
   gpc1_1 gpc1_1_1821(
      {stage38[96]},
      {stage38[109]}
   );
   gpc1_1 gpc1_1_1822(
      {stage38[97]},
      {stage38[110]}
   );
   gpc1_1 gpc1_1_1823(
      {stage38[98]},
      {stage38[111]}
   );
   gpc1_1 gpc1_1_1824(
      {stage38[99]},
      {stage38[112]}
   );
   gpc215_4 gpc215_4_1825(
      {stage38[100], stage38[101], stage38[102], stage38[103], stage38[104]},
      {stage39[94]},
      {stage40[101], stage40[102]},
      {stage41[127], stage40[122], stage39[106], stage38[113]}
   );
   gpc615_5 gpc615_5_1826(
      {stage39[95], stage39[96], stage39[97], stage39[98], stage39[99]},
      {stage40[103]},
      {stage41[110], stage41[111], stage41[112], stage41[113], stage41[114], stage41[115]},
      {stage43[128], stage42[130], stage41[128], stage40[123], stage39[107]}
   );
   gpc1406_5 gpc1406_5_1827(
      {stage39[100], stage39[101], stage39[102], stage39[103], 1'h0, 1'h0},
      {stage41[116], stage41[117], stage41[118], stage41[119]},
      {stage42[106]},
      {stage43[129], stage42[131], stage41[129], stage40[124], stage39[108]}
   );
   gpc1_1 gpc1_1_1828(
      {stage40[104]},
      {stage40[125]}
   );
   gpc1_1 gpc1_1_1829(
      {stage40[105]},
      {stage40[126]}
   );
   gpc1_1 gpc1_1_1830(
      {stage40[106]},
      {stage40[127]}
   );
   gpc1_1 gpc1_1_1831(
      {stage40[107]},
      {stage40[128]}
   );
   gpc606_5 gpc606_5_1832(
      {stage40[108], stage40[109], stage40[110], stage40[111], stage40[112], stage40[113]},
      {stage42[107], stage42[108], stage42[109], stage42[110], stage42[111], stage42[112]},
      {stage44[109], stage43[130], stage42[132], stage41[130], stage40[129]}
   );
   gpc606_5 gpc606_5_1833(
      {stage40[114], stage40[115], stage40[116], stage40[117], stage40[118], stage40[119]},
      {stage42[113], stage42[114], stage42[115], stage42[116], stage42[117], stage42[118]},
      {stage44[110], stage43[131], stage42[133], stage41[131], stage40[130]}
   );
   gpc1_1 gpc1_1_1834(
      {stage41[120]},
      {stage41[132]}
   );
   gpc1_1 gpc1_1_1835(
      {stage41[121]},
      {stage41[133]}
   );
   gpc1_1 gpc1_1_1836(
      {stage41[122]},
      {stage41[134]}
   );
   gpc1_1 gpc1_1_1837(
      {stage41[123]},
      {stage41[135]}
   );
   gpc1_1 gpc1_1_1838(
      {stage41[124]},
      {stage41[136]}
   );
   gpc1_1 gpc1_1_1839(
      {stage41[125]},
      {stage41[137]}
   );
   gpc1_1 gpc1_1_1840(
      {stage41[126]},
      {stage41[138]}
   );
   gpc1_1 gpc1_1_1841(
      {stage42[119]},
      {stage42[134]}
   );
   gpc615_5 gpc615_5_1842(
      {stage42[120], stage42[121], stage42[122], stage42[123], stage42[124]},
      {stage43[99]},
      {stage44[85], stage44[86], stage44[87], stage44[88], stage44[89], stage44[90]},
      {stage46[117], stage45[122], stage44[111], stage43[132], stage42[135]}
   );
   gpc615_5 gpc615_5_1843(
      {stage42[125], stage42[126], stage42[127], stage42[128], stage42[129]},
      {stage43[100]},
      {stage44[91], stage44[92], stage44[93], stage44[94], stage44[95], stage44[96]},
      {stage46[118], stage45[123], stage44[112], stage43[133], stage42[136]}
   );
   gpc1_1 gpc1_1_1844(
      {stage43[101]},
      {stage43[134]}
   );
   gpc1_1 gpc1_1_1845(
      {stage43[102]},
      {stage43[135]}
   );
   gpc1_1 gpc1_1_1846(
      {stage43[103]},
      {stage43[136]}
   );
   gpc1_1 gpc1_1_1847(
      {stage43[104]},
      {stage43[137]}
   );
   gpc1_1 gpc1_1_1848(
      {stage43[105]},
      {stage43[138]}
   );
   gpc1_1 gpc1_1_1849(
      {stage43[106]},
      {stage43[139]}
   );
   gpc1_1 gpc1_1_1850(
      {stage43[107]},
      {stage43[140]}
   );
   gpc1_1 gpc1_1_1851(
      {stage43[108]},
      {stage43[141]}
   );
   gpc1_1 gpc1_1_1852(
      {stage43[109]},
      {stage43[142]}
   );
   gpc1_1 gpc1_1_1853(
      {stage43[110]},
      {stage43[143]}
   );
   gpc1_1 gpc1_1_1854(
      {stage43[111]},
      {stage43[144]}
   );
   gpc1_1 gpc1_1_1855(
      {stage43[112]},
      {stage43[145]}
   );
   gpc1_1 gpc1_1_1856(
      {stage43[113]},
      {stage43[146]}
   );
   gpc1_1 gpc1_1_1857(
      {stage43[114]},
      {stage43[147]}
   );
   gpc1_1 gpc1_1_1858(
      {stage43[115]},
      {stage43[148]}
   );
   gpc606_5 gpc606_5_1859(
      {stage43[116], stage43[117], stage43[118], stage43[119], stage43[120], stage43[121]},
      {stage45[93], stage45[94], stage45[95], stage45[96], stage45[97], stage45[98]},
      {stage47[117], stage46[119], stage45[124], stage44[113], stage43[149]}
   );
   gpc606_5 gpc606_5_1860(
      {stage43[122], stage43[123], stage43[124], stage43[125], stage43[126], stage43[127]},
      {stage45[99], stage45[100], stage45[101], stage45[102], stage45[103], stage45[104]},
      {stage47[118], stage46[120], stage45[125], stage44[114], stage43[150]}
   );
   gpc606_5 gpc606_5_1861(
      {stage44[97], stage44[98], stage44[99], stage44[100], stage44[101], stage44[102]},
      {stage46[106], stage46[107], stage46[108], stage46[109], stage46[110], stage46[111]},
      {stage48[113], stage47[119], stage46[121], stage45[126], stage44[115]}
   );
   gpc606_5 gpc606_5_1862(
      {stage44[103], stage44[104], stage44[105], stage44[106], stage44[107], stage44[108]},
      {stage46[112], stage46[113], stage46[114], stage46[115], stage46[116], 1'h0},
      {stage48[114], stage47[120], stage46[122], stage45[127], stage44[116]}
   );
   gpc1_1 gpc1_1_1863(
      {stage45[105]},
      {stage45[128]}
   );
   gpc1_1 gpc1_1_1864(
      {stage45[106]},
      {stage45[129]}
   );
   gpc1_1 gpc1_1_1865(
      {stage45[107]},
      {stage45[130]}
   );
   gpc1_1 gpc1_1_1866(
      {stage45[108]},
      {stage45[131]}
   );
   gpc1_1 gpc1_1_1867(
      {stage45[109]},
      {stage45[132]}
   );
   gpc606_5 gpc606_5_1868(
      {stage45[110], stage45[111], stage45[112], stage45[113], stage45[114], stage45[115]},
      {stage47[91], stage47[92], stage47[93], stage47[94], stage47[95], stage47[96]},
      {stage49[117], stage48[115], stage47[121], stage46[123], stage45[133]}
   );
   gpc606_5 gpc606_5_1869(
      {stage45[116], stage45[117], stage45[118], stage45[119], stage45[120], stage45[121]},
      {stage47[97], stage47[98], stage47[99], stage47[100], stage47[101], stage47[102]},
      {stage49[118], stage48[116], stage47[122], stage46[124], stage45[134]}
   );
   gpc615_5 gpc615_5_1870(
      {stage47[103], stage47[104], stage47[105], stage47[106], stage47[107]},
      {stage48[101]},
      {stage49[89], stage49[90], stage49[91], stage49[92], stage49[93], stage49[94]},
      {stage51[103], stage50[110], stage49[119], stage48[117], stage47[123]}
   );
   gpc615_5 gpc615_5_1871(
      {stage47[108], stage47[109], stage47[110], stage47[111], stage47[112]},
      {stage48[102]},
      {stage49[95], stage49[96], stage49[97], stage49[98], stage49[99], stage49[100]},
      {stage51[104], stage50[111], stage49[120], stage48[118], stage47[124]}
   );
   gpc615_5 gpc615_5_1872(
      {stage47[113], stage47[114], stage47[115], stage47[116], 1'h0},
      {stage48[103]},
      {stage49[101], stage49[102], stage49[103], stage49[104], stage49[105], stage49[106]},
      {stage51[105], stage50[112], stage49[121], stage48[119], stage47[125]}
   );
   gpc1_1 gpc1_1_1873(
      {stage48[104]},
      {stage48[120]}
   );
   gpc1_1 gpc1_1_1874(
      {stage48[105]},
      {stage48[121]}
   );
   gpc1_1 gpc1_1_1875(
      {stage48[106]},
      {stage48[122]}
   );
   gpc606_5 gpc606_5_1876(
      {stage48[107], stage48[108], stage48[109], stage48[110], stage48[111], stage48[112]},
      {stage50[96], stage50[97], stage50[98], stage50[99], stage50[100], stage50[101]},
      {stage52[110], stage51[106], stage50[113], stage49[122], stage48[123]}
   );
   gpc1_1 gpc1_1_1877(
      {stage49[107]},
      {stage49[123]}
   );
   gpc1_1 gpc1_1_1878(
      {stage49[108]},
      {stage49[124]}
   );
   gpc1_1 gpc1_1_1879(
      {stage49[109]},
      {stage49[125]}
   );
   gpc1_1 gpc1_1_1880(
      {stage49[110]},
      {stage49[126]}
   );
   gpc1_1 gpc1_1_1881(
      {stage49[111]},
      {stage49[127]}
   );
   gpc1_1 gpc1_1_1882(
      {stage49[112]},
      {stage49[128]}
   );
   gpc1_1 gpc1_1_1883(
      {stage49[113]},
      {stage49[129]}
   );
   gpc1_1 gpc1_1_1884(
      {stage49[114]},
      {stage49[130]}
   );
   gpc1_1 gpc1_1_1885(
      {stage49[115]},
      {stage49[131]}
   );
   gpc1_1 gpc1_1_1886(
      {stage49[116]},
      {stage49[132]}
   );
   gpc615_5 gpc615_5_1887(
      {stage50[102], stage50[103], stage50[104], stage50[105], stage50[106]},
      {stage51[88]},
      {stage52[92], stage52[93], stage52[94], stage52[95], stage52[96], stage52[97]},
      {stage54[115], stage53[112], stage52[111], stage51[107], stage50[114]}
   );
   gpc615_5 gpc615_5_1888(
      {stage50[107], stage50[108], stage50[109], 1'h0, 1'h0},
      {stage51[89]},
      {stage52[98], stage52[99], stage52[100], stage52[101], stage52[102], stage52[103]},
      {stage54[116], stage53[113], stage52[112], stage51[108], stage50[115]}
   );
   gpc1_1 gpc1_1_1889(
      {stage51[90]},
      {stage51[109]}
   );
   gpc1_1 gpc1_1_1890(
      {stage51[91]},
      {stage51[110]}
   );
   gpc606_5 gpc606_5_1891(
      {stage51[92], stage51[93], stage51[94], stage51[95], stage51[96], stage51[97]},
      {stage53[95], stage53[96], stage53[97], stage53[98], stage53[99], stage53[100]},
      {stage55[107], stage54[117], stage53[114], stage52[113], stage51[111]}
   );
   gpc615_5 gpc615_5_1892(
      {stage51[98], stage51[99], stage51[100], stage51[101], stage51[102]},
      {stage52[104]},
      {stage53[101], stage53[102], stage53[103], stage53[104], stage53[105], stage53[106]},
      {stage55[108], stage54[118], stage53[115], stage52[114], stage51[112]}
   );
   gpc606_5 gpc606_5_1893(
      {stage52[105], stage52[106], stage52[107], stage52[108], stage52[109], 1'h0},
      {stage54[98], stage54[99], stage54[100], stage54[101], stage54[102], stage54[103]},
      {stage56[130], stage55[109], stage54[119], stage53[116], stage52[115]}
   );
   gpc135_4 gpc135_4_1894(
      {stage53[107], stage53[108], stage53[109], stage53[110], stage53[111]},
      {stage54[104], stage54[105], stage54[106]},
      {stage55[94]},
      {stage56[131], stage55[110], stage54[120], stage53[117]}
   );
   gpc1_1 gpc1_1_1895(
      {stage54[107]},
      {stage54[121]}
   );
   gpc1_1 gpc1_1_1896(
      {stage54[108]},
      {stage54[122]}
   );
   gpc1_1 gpc1_1_1897(
      {stage54[109]},
      {stage54[123]}
   );
   gpc615_5 gpc615_5_1898(
      {stage54[110], stage54[111], stage54[112], stage54[113], stage54[114]},
      {stage55[95]},
      {stage56[105], stage56[106], stage56[107], stage56[108], stage56[109], stage56[110]},
      {stage58[114], stage57[108], stage56[132], stage55[111], stage54[124]}
   );
   gpc606_5 gpc606_5_1899(
      {stage55[96], stage55[97], stage55[98], stage55[99], stage55[100], stage55[101]},
      {stage57[92], stage57[93], stage57[94], stage57[95], stage57[96], stage57[97]},
      {stage59[121], stage58[115], stage57[109], stage56[133], stage55[112]}
   );
   gpc606_5 gpc606_5_1900(
      {stage55[102], stage55[103], stage55[104], stage55[105], stage55[106], 1'h0},
      {stage57[98], stage57[99], stage57[100], stage57[101], stage57[102], stage57[103]},
      {stage59[122], stage58[116], stage57[110], stage56[134], stage55[113]}
   );
   gpc1_1 gpc1_1_1901(
      {stage56[111]},
      {stage56[135]}
   );
   gpc1_1 gpc1_1_1902(
      {stage56[112]},
      {stage56[136]}
   );
   gpc1_1 gpc1_1_1903(
      {stage56[113]},
      {stage56[137]}
   );
   gpc1_1 gpc1_1_1904(
      {stage56[114]},
      {stage56[138]}
   );
   gpc1_1 gpc1_1_1905(
      {stage56[115]},
      {stage56[139]}
   );
   gpc1_1 gpc1_1_1906(
      {stage56[116]},
      {stage56[140]}
   );
   gpc1_1 gpc1_1_1907(
      {stage56[117]},
      {stage56[141]}
   );
   gpc1_1 gpc1_1_1908(
      {stage56[118]},
      {stage56[142]}
   );
   gpc1_1 gpc1_1_1909(
      {stage56[119]},
      {stage56[143]}
   );
   gpc615_5 gpc615_5_1910(
      {stage56[120], stage56[121], stage56[122], stage56[123], stage56[124]},
      {stage57[104]},
      {stage58[99], stage58[100], stage58[101], stage58[102], stage58[103], stage58[104]},
      {stage60[117], stage59[123], stage58[117], stage57[111], stage56[144]}
   );
   gpc615_5 gpc615_5_1911(
      {stage56[125], stage56[126], stage56[127], stage56[128], stage56[129]},
      {stage57[105]},
      {stage58[105], stage58[106], stage58[107], stage58[108], stage58[109], stage58[110]},
      {stage60[118], stage59[124], stage58[118], stage57[112], stage56[145]}
   );
   gpc606_5 gpc606_5_1912(
      {stage57[106], stage57[107], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage59[99], stage59[100], stage59[101], stage59[102], stage59[103], stage59[104]},
      {stage61[125], stage60[119], stage59[125], stage58[119], stage57[113]}
   );
   gpc615_5 gpc615_5_1913(
      {stage58[111], stage58[112], stage58[113], 1'h0, 1'h0},
      {stage59[105]},
      {stage60[98], stage60[99], stage60[100], stage60[101], stage60[102], stage60[103]},
      {stage62[110], stage61[126], stage60[120], stage59[126], stage58[120]}
   );
   gpc606_5 gpc606_5_1914(
      {stage59[106], stage59[107], stage59[108], stage59[109], stage59[110], stage59[111]},
      {stage61[104], stage61[105], stage61[106], stage61[107], stage61[108], stage61[109]},
      {stage63[110], stage62[111], stage61[127], stage60[121], stage59[127]}
   );
   gpc135_4 gpc135_4_1915(
      {stage59[112], stage59[113], stage59[114], stage59[115], stage59[116]},
      {stage60[104], stage60[105], stage60[106]},
      {stage61[110]},
      {stage62[112], stage61[128], stage60[122], stage59[128]}
   );
   gpc135_4 gpc135_4_1916(
      {stage59[117], stage59[118], stage59[119], stage59[120], 1'h0},
      {stage60[107], stage60[108], stage60[109]},
      {stage61[111]},
      {stage62[113], stage61[129], stage60[123], stage59[129]}
   );
   gpc1_1 gpc1_1_1917(
      {stage60[110]},
      {stage60[124]}
   );
   gpc1_1 gpc1_1_1918(
      {stage60[111]},
      {stage60[125]}
   );
   gpc1_1 gpc1_1_1919(
      {stage60[112]},
      {stage60[126]}
   );
   gpc1_1 gpc1_1_1920(
      {stage60[113]},
      {stage60[127]}
   );
   gpc1_1 gpc1_1_1921(
      {stage60[114]},
      {stage60[128]}
   );
   gpc1_1 gpc1_1_1922(
      {stage60[115]},
      {stage60[129]}
   );
   gpc1_1 gpc1_1_1923(
      {stage60[116]},
      {stage60[130]}
   );
   gpc1_1 gpc1_1_1924(
      {stage61[112]},
      {stage61[130]}
   );
   gpc606_5 gpc606_5_1925(
      {stage61[113], stage61[114], stage61[115], stage61[116], stage61[117], stage61[118]},
      {stage63[97], stage63[98], stage63[99], stage63[100], stage63[101], stage63[102]},
      {stage65[16], stage64[31], stage63[111], stage62[114], stage61[131]}
   );
   gpc606_5 gpc606_5_1926(
      {stage61[119], stage61[120], stage61[121], stage61[122], stage61[123], stage61[124]},
      {stage63[103], stage63[104], stage63[105], stage63[106], stage63[107], stage63[108]},
      {stage65[17], stage64[32], stage63[112], stage62[115], stage61[132]}
   );
   gpc1_1 gpc1_1_1927(
      {stage62[93]},
      {stage62[116]}
   );
   gpc1_1 gpc1_1_1928(
      {stage62[94]},
      {stage62[117]}
   );
   gpc1_1 gpc1_1_1929(
      {stage62[95]},
      {stage62[118]}
   );
   gpc1_1 gpc1_1_1930(
      {stage62[96]},
      {stage62[119]}
   );
   gpc1_1 gpc1_1_1931(
      {stage62[97]},
      {stage62[120]}
   );
   gpc1_1 gpc1_1_1932(
      {stage62[98]},
      {stage62[121]}
   );
   gpc1_1 gpc1_1_1933(
      {stage62[99]},
      {stage62[122]}
   );
   gpc1_1 gpc1_1_1934(
      {stage62[100]},
      {stage62[123]}
   );
   gpc1_1 gpc1_1_1935(
      {stage62[101]},
      {stage62[124]}
   );
   gpc1_1 gpc1_1_1936(
      {stage62[102]},
      {stage62[125]}
   );
   gpc1_1 gpc1_1_1937(
      {stage62[103]},
      {stage62[126]}
   );
   gpc606_5 gpc606_5_1938(
      {stage62[104], stage62[105], stage62[106], stage62[107], stage62[108], stage62[109]},
      {stage64[16], stage64[17], stage64[18], stage64[19], stage64[20], stage64[21]},
      {stage66[3], stage65[18], stage64[33], stage63[113], stage62[127]}
   );
   gpc1_1 gpc1_1_1939(
      {stage63[109]},
      {stage63[114]}
   );
   gpc1_1 gpc1_1_1940(
      {stage64[22]},
      {stage64[34]}
   );
   gpc1_1 gpc1_1_1941(
      {stage64[23]},
      {stage64[35]}
   );
   gpc1_1 gpc1_1_1942(
      {stage64[24]},
      {stage64[36]}
   );
   gpc1_1 gpc1_1_1943(
      {stage64[25]},
      {stage64[37]}
   );
   gpc1_1 gpc1_1_1944(
      {stage64[26]},
      {stage64[38]}
   );
   gpc1_1 gpc1_1_1945(
      {stage64[27]},
      {stage64[39]}
   );
   gpc1_1 gpc1_1_1946(
      {stage64[28]},
      {stage64[40]}
   );
   gpc1_1 gpc1_1_1947(
      {stage64[29]},
      {stage64[41]}
   );
   gpc1_1 gpc1_1_1948(
      {stage64[30]},
      {stage64[42]}
   );
   gpc1_1 gpc1_1_1949(
      {stage65[8]},
      {stage65[19]}
   );
   gpc1_1 gpc1_1_1950(
      {stage65[9]},
      {stage65[20]}
   );
   gpc1_1 gpc1_1_1951(
      {stage65[10]},
      {stage65[21]}
   );
   gpc1_1 gpc1_1_1952(
      {stage65[11]},
      {stage65[22]}
   );
   gpc1_1 gpc1_1_1953(
      {stage65[12]},
      {stage65[23]}
   );
   gpc1_1 gpc1_1_1954(
      {stage65[13]},
      {stage65[24]}
   );
   gpc1_1 gpc1_1_1955(
      {stage65[14]},
      {stage65[25]}
   );
   gpc1_1 gpc1_1_1956(
      {stage65[15]},
      {stage65[26]}
   );
   gpc1_1 gpc1_1_1957(
      {stage66[0]},
      {stage66[4]}
   );
   gpc1_1 gpc1_1_1958(
      {stage66[1]},
      {stage66[5]}
   );
   gpc1_1 gpc1_1_1959(
      {stage66[2]},
      {stage66[6]}
   );
   gpc1_1 gpc1_1_1960(
      {stage67[0]},
      {stage67[1]}
   );
   gpc1_1 gpc1_1_1961(
      {stage00[86]},
      {stage00[92]}
   );
   gpc1_1 gpc1_1_1962(
      {stage00[87]},
      {stage00[93]}
   );
   gpc1_1 gpc1_1_1963(
      {stage00[88]},
      {stage00[94]}
   );
   gpc1_1 gpc1_1_1964(
      {stage00[89]},
      {stage00[95]}
   );
   gpc1_1 gpc1_1_1965(
      {stage00[90]},
      {stage00[96]}
   );
   gpc1_1 gpc1_1_1966(
      {stage00[91]},
      {stage00[97]}
   );
   gpc1_1 gpc1_1_1967(
      {stage01[123]},
      {stage01[126]}
   );
   gpc1_1 gpc1_1_1968(
      {stage01[124]},
      {stage01[127]}
   );
   gpc1_1 gpc1_1_1969(
      {stage01[125]},
      {stage01[128]}
   );
   gpc1_1 gpc1_1_1970(
      {stage02[105]},
      {stage02[111]}
   );
   gpc1_1 gpc1_1_1971(
      {stage02[106]},
      {stage02[112]}
   );
   gpc1_1 gpc1_1_1972(
      {stage02[107]},
      {stage02[113]}
   );
   gpc1_1 gpc1_1_1973(
      {stage02[108]},
      {stage02[114]}
   );
   gpc1_1 gpc1_1_1974(
      {stage02[109]},
      {stage02[115]}
   );
   gpc1_1 gpc1_1_1975(
      {stage02[110]},
      {stage02[116]}
   );
   gpc615_5 gpc615_5_1976(
      {stage03[133], stage03[134], stage03[135], stage03[136], stage03[137]},
      {stage04[112]},
      {stage05[111], stage05[112], stage05[113], stage05[114], stage05[115], stage05[116]},
      {stage07[115], stage06[109], stage05[122], stage04[118], stage03[138]}
   );
   gpc1_1 gpc1_1_1977(
      {stage04[113]},
      {stage04[119]}
   );
   gpc1_1 gpc1_1_1978(
      {stage04[114]},
      {stage04[120]}
   );
   gpc1_1 gpc1_1_1979(
      {stage04[115]},
      {stage04[121]}
   );
   gpc1_1 gpc1_1_1980(
      {stage04[116]},
      {stage04[122]}
   );
   gpc1_1 gpc1_1_1981(
      {stage04[117]},
      {stage04[123]}
   );
   gpc1_1 gpc1_1_1982(
      {stage05[117]},
      {stage05[123]}
   );
   gpc1_1 gpc1_1_1983(
      {stage05[118]},
      {stage05[124]}
   );
   gpc1_1 gpc1_1_1984(
      {stage05[119]},
      {stage05[125]}
   );
   gpc1_1 gpc1_1_1985(
      {stage05[120]},
      {stage05[126]}
   );
   gpc1_1 gpc1_1_1986(
      {stage05[121]},
      {stage05[127]}
   );
   gpc1_1 gpc1_1_1987(
      {stage06[99]},
      {stage06[110]}
   );
   gpc1_1 gpc1_1_1988(
      {stage06[100]},
      {stage06[111]}
   );
   gpc1_1 gpc1_1_1989(
      {stage06[101]},
      {stage06[112]}
   );
   gpc7_3 gpc7_3_1990(
      {stage06[102], stage06[103], stage06[104], stage06[105], stage06[106], stage06[107], stage06[108]},
      {stage08[125], stage07[116], stage06[113]}
   );
   gpc1_1 gpc1_1_1991(
      {stage07[111]},
      {stage07[117]}
   );
   gpc1_1 gpc1_1_1992(
      {stage07[112]},
      {stage07[118]}
   );
   gpc1_1 gpc1_1_1993(
      {stage07[113]},
      {stage07[119]}
   );
   gpc1_1 gpc1_1_1994(
      {stage07[114]},
      {stage07[120]}
   );
   gpc606_5 gpc606_5_1995(
      {stage08[119], stage08[120], stage08[121], stage08[122], stage08[123], stage08[124]},
      {stage10[130], stage10[131], stage10[132], stage10[133], stage10[134], stage10[135]},
      {stage12[143], stage11[153], stage10[139], stage09[167], stage08[126]}
   );
   gpc1_1 gpc1_1_1996(
      {stage09[152]},
      {stage09[168]}
   );
   gpc1_1 gpc1_1_1997(
      {stage09[153]},
      {stage09[169]}
   );
   gpc1_1 gpc1_1_1998(
      {stage09[154]},
      {stage09[170]}
   );
   gpc606_5 gpc606_5_1999(
      {stage09[155], stage09[156], stage09[157], stage09[158], stage09[159], stage09[160]},
      {stage11[134], stage11[135], stage11[136], stage11[137], stage11[138], stage11[139]},
      {stage13[126], stage12[144], stage11[154], stage10[140], stage09[171]}
   );
   gpc606_5 gpc606_5_2000(
      {stage09[161], stage09[162], stage09[163], stage09[164], stage09[165], stage09[166]},
      {stage11[140], stage11[141], stage11[142], stage11[143], stage11[144], stage11[145]},
      {stage13[127], stage12[145], stage11[155], stage10[141], stage09[172]}
   );
   gpc1_1 gpc1_1_2001(
      {stage10[136]},
      {stage10[142]}
   );
   gpc1_1 gpc1_1_2002(
      {stage10[137]},
      {stage10[143]}
   );
   gpc1_1 gpc1_1_2003(
      {stage10[138]},
      {stage10[144]}
   );
   gpc1_1 gpc1_1_2004(
      {stage11[146]},
      {stage11[156]}
   );
   gpc606_5 gpc606_5_2005(
      {stage11[147], stage11[148], stage11[149], stage11[150], stage11[151], stage11[152]},
      {stage13[107], stage13[108], stage13[109], stage13[110], stage13[111], stage13[112]},
      {stage15[156], stage14[110], stage13[128], stage12[146], stage11[157]}
   );
   gpc1_1 gpc1_1_2006(
      {stage12[131]},
      {stage12[147]}
   );
   gpc1_1 gpc1_1_2007(
      {stage12[132]},
      {stage12[148]}
   );
   gpc135_4 gpc135_4_2008(
      {stage12[133], stage12[134], stage12[135], stage12[136], stage12[137]},
      {stage13[113], stage13[114], stage13[115]},
      {stage14[105]},
      {stage15[157], stage14[111], stage13[129], stage12[149]}
   );
   gpc135_4 gpc135_4_2009(
      {stage12[138], stage12[139], stage12[140], stage12[141], stage12[142]},
      {stage13[116], stage13[117], stage13[118]},
      {stage14[106]},
      {stage15[158], stage14[112], stage13[130], stage12[150]}
   );
   gpc1_1 gpc1_1_2010(
      {stage13[119]},
      {stage13[131]}
   );
   gpc1_1 gpc1_1_2011(
      {stage13[120]},
      {stage13[132]}
   );
   gpc1_1 gpc1_1_2012(
      {stage13[121]},
      {stage13[133]}
   );
   gpc1_1 gpc1_1_2013(
      {stage13[122]},
      {stage13[134]}
   );
   gpc1_1 gpc1_1_2014(
      {stage13[123]},
      {stage13[135]}
   );
   gpc1_1 gpc1_1_2015(
      {stage13[124]},
      {stage13[136]}
   );
   gpc1_1 gpc1_1_2016(
      {stage13[125]},
      {stage13[137]}
   );
   gpc1_1 gpc1_1_2017(
      {stage14[107]},
      {stage14[113]}
   );
   gpc1_1 gpc1_1_2018(
      {stage14[108]},
      {stage14[114]}
   );
   gpc1_1 gpc1_1_2019(
      {stage14[109]},
      {stage14[115]}
   );
   gpc1_1 gpc1_1_2020(
      {stage15[145]},
      {stage15[159]}
   );
   gpc1_1 gpc1_1_2021(
      {stage15[146]},
      {stage15[160]}
   );
   gpc1_1 gpc1_1_2022(
      {stage15[147]},
      {stage15[161]}
   );
   gpc1_1 gpc1_1_2023(
      {stage15[148]},
      {stage15[162]}
   );
   gpc1_1 gpc1_1_2024(
      {stage15[149]},
      {stage15[163]}
   );
   gpc1_1 gpc1_1_2025(
      {stage15[150]},
      {stage15[164]}
   );
   gpc615_5 gpc615_5_2026(
      {stage15[151], stage15[152], stage15[153], stage15[154], stage15[155]},
      {stage16[105]},
      {stage17[138], stage17[139], stage17[140], stage17[141], stage17[142], stage17[143]},
      {stage19[122], stage18[120], stage17[149], stage16[111], stage15[165]}
   );
   gpc135_4 gpc135_4_2027(
      {stage16[106], stage16[107], stage16[108], stage16[109], stage16[110]},
      {stage17[144], stage17[145], stage17[146]},
      {stage18[102]},
      {stage19[123], stage18[121], stage17[150], stage16[112]}
   );
   gpc1_1 gpc1_1_2028(
      {stage17[147]},
      {stage17[151]}
   );
   gpc1_1 gpc1_1_2029(
      {stage17[148]},
      {stage17[152]}
   );
   gpc1_1 gpc1_1_2030(
      {stage18[103]},
      {stage18[122]}
   );
   gpc1_1 gpc1_1_2031(
      {stage18[104]},
      {stage18[123]}
   );
   gpc615_5 gpc615_5_2032(
      {stage18[105], stage18[106], stage18[107], stage18[108], stage18[109]},
      {stage19[115]},
      {stage20[125], stage20[126], stage20[127], stage20[128], stage20[129], stage20[130]},
      {stage22[113], stage21[112], stage20[147], stage19[124], stage18[124]}
   );
   gpc615_5 gpc615_5_2033(
      {stage18[110], stage18[111], stage18[112], stage18[113], stage18[114]},
      {stage19[116]},
      {stage20[131], stage20[132], stage20[133], stage20[134], stage20[135], stage20[136]},
      {stage22[114], stage21[113], stage20[148], stage19[125], stage18[125]}
   );
   gpc615_5 gpc615_5_2034(
      {stage18[115], stage18[116], stage18[117], stage18[118], stage18[119]},
      {stage19[117]},
      {stage20[137], stage20[138], stage20[139], stage20[140], stage20[141], stage20[142]},
      {stage22[115], stage21[114], stage20[149], stage19[126], stage18[126]}
   );
   gpc1_1 gpc1_1_2035(
      {stage19[118]},
      {stage19[127]}
   );
   gpc1_1 gpc1_1_2036(
      {stage19[119]},
      {stage19[128]}
   );
   gpc1_1 gpc1_1_2037(
      {stage19[120]},
      {stage19[129]}
   );
   gpc1_1 gpc1_1_2038(
      {stage19[121]},
      {stage19[130]}
   );
   gpc1_1 gpc1_1_2039(
      {stage20[143]},
      {stage20[150]}
   );
   gpc1_1 gpc1_1_2040(
      {stage20[144]},
      {stage20[151]}
   );
   gpc1_1 gpc1_1_2041(
      {stage20[145]},
      {stage20[152]}
   );
   gpc1_1 gpc1_1_2042(
      {stage20[146]},
      {stage20[153]}
   );
   gpc1_1 gpc1_1_2043(
      {stage21[105]},
      {stage21[115]}
   );
   gpc1_1 gpc1_1_2044(
      {stage21[106]},
      {stage21[116]}
   );
   gpc215_4 gpc215_4_2045(
      {stage21[107], stage21[108], stage21[109], stage21[110], stage21[111]},
      {stage22[109]},
      {stage23[119], stage23[120]},
      {stage24[117], stage23[135], stage22[116], stage21[117]}
   );
   gpc1_1 gpc1_1_2046(
      {stage22[110]},
      {stage22[117]}
   );
   gpc1_1 gpc1_1_2047(
      {stage22[111]},
      {stage22[118]}
   );
   gpc1_1 gpc1_1_2048(
      {stage22[112]},
      {stage22[119]}
   );
   gpc1_1 gpc1_1_2049(
      {stage23[121]},
      {stage23[136]}
   );
   gpc1_1 gpc1_1_2050(
      {stage23[122]},
      {stage23[137]}
   );
   gpc1_1 gpc1_1_2051(
      {stage23[123]},
      {stage23[138]}
   );
   gpc606_5 gpc606_5_2052(
      {stage23[124], stage23[125], stage23[126], stage23[127], stage23[128], stage23[129]},
      {stage25[117], stage25[118], stage25[119], stage25[120], stage25[121], stage25[122]},
      {stage27[136], stage26[103], stage25[132], stage24[118], stage23[139]}
   );
   gpc615_5 gpc615_5_2053(
      {stage23[130], stage23[131], stage23[132], stage23[133], stage23[134]},
      {stage24[112]},
      {stage25[123], stage25[124], stage25[125], stage25[126], stage25[127], stage25[128]},
      {stage27[137], stage26[104], stage25[133], stage24[119], stage23[140]}
   );
   gpc1_1 gpc1_1_2054(
      {stage24[113]},
      {stage24[120]}
   );
   gpc1_1 gpc1_1_2055(
      {stage24[114]},
      {stage24[121]}
   );
   gpc1_1 gpc1_1_2056(
      {stage24[115]},
      {stage24[122]}
   );
   gpc1_1 gpc1_1_2057(
      {stage24[116]},
      {stage24[123]}
   );
   gpc1_1 gpc1_1_2058(
      {stage25[129]},
      {stage25[134]}
   );
   gpc1_1 gpc1_1_2059(
      {stage25[130]},
      {stage25[135]}
   );
   gpc1_1 gpc1_1_2060(
      {stage25[131]},
      {stage25[136]}
   );
   gpc1_1 gpc1_1_2061(
      {stage26[96]},
      {stage26[105]}
   );
   gpc1_1 gpc1_1_2062(
      {stage26[97]},
      {stage26[106]}
   );
   gpc1_1 gpc1_1_2063(
      {stage26[98]},
      {stage26[107]}
   );
   gpc1_1 gpc1_1_2064(
      {stage26[99]},
      {stage26[108]}
   );
   gpc1_1 gpc1_1_2065(
      {stage26[100]},
      {stage26[109]}
   );
   gpc1_1 gpc1_1_2066(
      {stage26[101]},
      {stage26[110]}
   );
   gpc1_1 gpc1_1_2067(
      {stage26[102]},
      {stage26[111]}
   );
   gpc1_1 gpc1_1_2068(
      {stage27[127]},
      {stage27[138]}
   );
   gpc1_1 gpc1_1_2069(
      {stage27[128]},
      {stage27[139]}
   );
   gpc1_1 gpc1_1_2070(
      {stage27[129]},
      {stage27[140]}
   );
   gpc1_1 gpc1_1_2071(
      {stage27[130]},
      {stage27[141]}
   );
   gpc1_1 gpc1_1_2072(
      {stage27[131]},
      {stage27[142]}
   );
   gpc1_1 gpc1_1_2073(
      {stage27[132]},
      {stage27[143]}
   );
   gpc1_1 gpc1_1_2074(
      {stage27[133]},
      {stage27[144]}
   );
   gpc1_1 gpc1_1_2075(
      {stage27[134]},
      {stage27[145]}
   );
   gpc1_1 gpc1_1_2076(
      {stage27[135]},
      {stage27[146]}
   );
   gpc1_1 gpc1_1_2077(
      {stage28[125]},
      {stage28[138]}
   );
   gpc1_1 gpc1_1_2078(
      {stage28[126]},
      {stage28[139]}
   );
   gpc1_1 gpc1_1_2079(
      {stage28[127]},
      {stage28[140]}
   );
   gpc1_1 gpc1_1_2080(
      {stage28[128]},
      {stage28[141]}
   );
   gpc1_1 gpc1_1_2081(
      {stage28[129]},
      {stage28[142]}
   );
   gpc1_1 gpc1_1_2082(
      {stage28[130]},
      {stage28[143]}
   );
   gpc7_3 gpc7_3_2083(
      {stage28[131], stage28[132], stage28[133], stage28[134], stage28[135], stage28[136], stage28[137]},
      {stage30[129], stage29[107], stage28[144]}
   );
   gpc1_1 gpc1_1_2084(
      {stage29[99]},
      {stage29[108]}
   );
   gpc1_1 gpc1_1_2085(
      {stage29[100]},
      {stage29[109]}
   );
   gpc1_1 gpc1_1_2086(
      {stage29[101]},
      {stage29[110]}
   );
   gpc1_1 gpc1_1_2087(
      {stage29[102]},
      {stage29[111]}
   );
   gpc1_1 gpc1_1_2088(
      {stage29[103]},
      {stage29[112]}
   );
   gpc623_5 gpc623_5_2089(
      {stage29[104], stage29[105], stage29[106]},
      {stage30[121], stage30[122]},
      {stage31[107], stage31[108], stage31[109], stage31[110], stage31[111], stage31[112]},
      {stage33[110], stage32[111], stage31[122], stage30[130], stage29[113]}
   );
   gpc1_1 gpc1_1_2090(
      {stage30[123]},
      {stage30[131]}
   );
   gpc1_1 gpc1_1_2091(
      {stage30[124]},
      {stage30[132]}
   );
   gpc1_1 gpc1_1_2092(
      {stage30[125]},
      {stage30[133]}
   );
   gpc623_5 gpc623_5_2093(
      {stage30[126], stage30[127], stage30[128]},
      {stage31[113], stage31[114]},
      {stage32[105], stage32[106], stage32[107], stage32[108], stage32[109], stage32[110]},
      {stage34[109], stage33[111], stage32[112], stage31[123], stage30[134]}
   );
   gpc1_1 gpc1_1_2094(
      {stage31[115]},
      {stage31[124]}
   );
   gpc1406_5 gpc1406_5_2095(
      {stage31[116], stage31[117], stage31[118], stage31[119], stage31[120], stage31[121]},
      {stage33[106], stage33[107], stage33[108], stage33[109]},
      {stage34[102]},
      {stage35[112], stage34[110], stage33[112], stage32[113], stage31[125]}
   );
   gpc1_1 gpc1_1_2096(
      {stage34[103]},
      {stage34[111]}
   );
   gpc1_1 gpc1_1_2097(
      {stage34[104]},
      {stage34[112]}
   );
   gpc1_1 gpc1_1_2098(
      {stage34[105]},
      {stage34[113]}
   );
   gpc1_1 gpc1_1_2099(
      {stage34[106]},
      {stage34[114]}
   );
   gpc1_1 gpc1_1_2100(
      {stage34[107]},
      {stage34[115]}
   );
   gpc1_1 gpc1_1_2101(
      {stage34[108]},
      {stage34[116]}
   );
   gpc1_1 gpc1_1_2102(
      {stage35[106]},
      {stage35[113]}
   );
   gpc615_5 gpc615_5_2103(
      {stage35[107], stage35[108], stage35[109], stage35[110], stage35[111]},
      {stage36[121]},
      {stage37[109], stage37[110], stage37[111], stage37[112], stage37[113], stage37[114]},
      {stage39[109], stage38[114], stage37[120], stage36[132], stage35[114]}
   );
   gpc1_1 gpc1_1_2104(
      {stage36[122]},
      {stage36[133]}
   );
   gpc1_1 gpc1_1_2105(
      {stage36[123]},
      {stage36[134]}
   );
   gpc1_1 gpc1_1_2106(
      {stage36[124]},
      {stage36[135]}
   );
   gpc1_1 gpc1_1_2107(
      {stage36[125]},
      {stage36[136]}
   );
   gpc1_1 gpc1_1_2108(
      {stage36[126]},
      {stage36[137]}
   );
   gpc1_1 gpc1_1_2109(
      {stage36[127]},
      {stage36[138]}
   );
   gpc1_1 gpc1_1_2110(
      {stage36[128]},
      {stage36[139]}
   );
   gpc1_1 gpc1_1_2111(
      {stage36[129]},
      {stage36[140]}
   );
   gpc1_1 gpc1_1_2112(
      {stage36[130]},
      {stage36[141]}
   );
   gpc1_1 gpc1_1_2113(
      {stage36[131]},
      {stage36[142]}
   );
   gpc1_1 gpc1_1_2114(
      {stage37[115]},
      {stage37[121]}
   );
   gpc1_1 gpc1_1_2115(
      {stage37[116]},
      {stage37[122]}
   );
   gpc1_1 gpc1_1_2116(
      {stage37[117]},
      {stage37[123]}
   );
   gpc1_1 gpc1_1_2117(
      {stage37[118]},
      {stage37[124]}
   );
   gpc1_1 gpc1_1_2118(
      {stage37[119]},
      {stage37[125]}
   );
   gpc1_1 gpc1_1_2119(
      {stage38[105]},
      {stage38[115]}
   );
   gpc1_1 gpc1_1_2120(
      {stage38[106]},
      {stage38[116]}
   );
   gpc1_1 gpc1_1_2121(
      {stage38[107]},
      {stage38[117]}
   );
   gpc606_5 gpc606_5_2122(
      {stage38[108], stage38[109], stage38[110], stage38[111], stage38[112], stage38[113]},
      {stage40[120], stage40[121], stage40[122], stage40[123], stage40[124], stage40[125]},
      {stage42[137], stage41[139], stage40[131], stage39[110], stage38[118]}
   );
   gpc1_1 gpc1_1_2123(
      {stage39[104]},
      {stage39[111]}
   );
   gpc1_1 gpc1_1_2124(
      {stage39[105]},
      {stage39[112]}
   );
   gpc1_1 gpc1_1_2125(
      {stage39[106]},
      {stage39[113]}
   );
   gpc1_1 gpc1_1_2126(
      {stage39[107]},
      {stage39[114]}
   );
   gpc1_1 gpc1_1_2127(
      {stage39[108]},
      {stage39[115]}
   );
   gpc1_1 gpc1_1_2128(
      {stage40[126]},
      {stage40[132]}
   );
   gpc1_1 gpc1_1_2129(
      {stage40[127]},
      {stage40[133]}
   );
   gpc1_1 gpc1_1_2130(
      {stage40[128]},
      {stage40[134]}
   );
   gpc1_1 gpc1_1_2131(
      {stage40[129]},
      {stage40[135]}
   );
   gpc1_1 gpc1_1_2132(
      {stage40[130]},
      {stage40[136]}
   );
   gpc1_1 gpc1_1_2133(
      {stage41[127]},
      {stage41[140]}
   );
   gpc1_1 gpc1_1_2134(
      {stage41[128]},
      {stage41[141]}
   );
   gpc615_5 gpc615_5_2135(
      {stage41[129], stage41[130], stage41[131], stage41[132], stage41[133]},
      {stage42[130]},
      {stage43[128], stage43[129], stage43[130], stage43[131], stage43[132], stage43[133]},
      {stage45[135], stage44[117], stage43[151], stage42[138], stage41[142]}
   );
   gpc615_5 gpc615_5_2136(
      {stage41[134], stage41[135], stage41[136], stage41[137], stage41[138]},
      {stage42[131]},
      {stage43[134], stage43[135], stage43[136], stage43[137], stage43[138], stage43[139]},
      {stage45[136], stage44[118], stage43[152], stage42[139], stage41[143]}
   );
   gpc606_5 gpc606_5_2137(
      {stage42[132], stage42[133], stage42[134], stage42[135], stage42[136], 1'h0},
      {stage44[109], stage44[110], stage44[111], stage44[112], stage44[113], stage44[114]},
      {stage46[125], stage45[137], stage44[119], stage43[153], stage42[140]}
   );
   gpc1_1 gpc1_1_2138(
      {stage43[140]},
      {stage43[154]}
   );
   gpc615_5 gpc615_5_2139(
      {stage43[141], stage43[142], stage43[143], stage43[144], stage43[145]},
      {stage44[115]},
      {stage45[122], stage45[123], stage45[124], stage45[125], stage45[126], stage45[127]},
      {stage47[126], stage46[126], stage45[138], stage44[120], stage43[155]}
   );
   gpc615_5 gpc615_5_2140(
      {stage43[146], stage43[147], stage43[148], stage43[149], stage43[150]},
      {stage44[116]},
      {stage45[128], stage45[129], stage45[130], stage45[131], stage45[132], stage45[133]},
      {stage47[127], stage46[127], stage45[139], stage44[121], stage43[156]}
   );
   gpc1_1 gpc1_1_2141(
      {stage45[134]},
      {stage45[140]}
   );
   gpc615_5 gpc615_5_2142(
      {stage46[117], stage46[118], stage46[119], stage46[120], stage46[121]},
      {stage47[117]},
      {stage48[113], stage48[114], stage48[115], stage48[116], stage48[117], stage48[118]},
      {stage50[116], stage49[133], stage48[124], stage47[128], stage46[128]}
   );
   gpc1343_5 gpc1343_5_2143(
      {stage46[122], stage46[123], stage46[124]},
      {stage47[118], stage47[119], stage47[120], stage47[121]},
      {stage48[119], stage48[120], stage48[121]},
      {stage49[117]},
      {stage50[117], stage49[134], stage48[125], stage47[129], stage46[129]}
   );
   gpc1_1 gpc1_1_2144(
      {stage47[122]},
      {stage47[130]}
   );
   gpc1_1 gpc1_1_2145(
      {stage47[123]},
      {stage47[131]}
   );
   gpc1_1 gpc1_1_2146(
      {stage47[124]},
      {stage47[132]}
   );
   gpc1_1 gpc1_1_2147(
      {stage47[125]},
      {stage47[133]}
   );
   gpc1_1 gpc1_1_2148(
      {stage48[122]},
      {stage48[126]}
   );
   gpc1_1 gpc1_1_2149(
      {stage48[123]},
      {stage48[127]}
   );
   gpc1_1 gpc1_1_2150(
      {stage49[118]},
      {stage49[135]}
   );
   gpc1_1 gpc1_1_2151(
      {stage49[119]},
      {stage49[136]}
   );
   gpc1_1 gpc1_1_2152(
      {stage49[120]},
      {stage49[137]}
   );
   gpc1_1 gpc1_1_2153(
      {stage49[121]},
      {stage49[138]}
   );
   gpc1_1 gpc1_1_2154(
      {stage49[122]},
      {stage49[139]}
   );
   gpc1_1 gpc1_1_2155(
      {stage49[123]},
      {stage49[140]}
   );
   gpc1_1 gpc1_1_2156(
      {stage49[124]},
      {stage49[141]}
   );
   gpc1_1 gpc1_1_2157(
      {stage49[125]},
      {stage49[142]}
   );
   gpc1_1 gpc1_1_2158(
      {stage49[126]},
      {stage49[143]}
   );
   gpc606_5 gpc606_5_2159(
      {stage49[127], stage49[128], stage49[129], stage49[130], stage49[131], stage49[132]},
      {stage51[103], stage51[104], stage51[105], stage51[106], stage51[107], stage51[108]},
      {stage53[118], stage52[116], stage51[113], stage50[118], stage49[144]}
   );
   gpc1_1 gpc1_1_2160(
      {stage50[110]},
      {stage50[119]}
   );
   gpc615_5 gpc615_5_2161(
      {stage50[111], stage50[112], stage50[113], stage50[114], stage50[115]},
      {stage51[109]},
      {stage52[110], stage52[111], stage52[112], stage52[113], stage52[114], stage52[115]},
      {stage54[125], stage53[119], stage52[117], stage51[114], stage50[120]}
   );
   gpc1_1 gpc1_1_2162(
      {stage51[110]},
      {stage51[115]}
   );
   gpc1_1 gpc1_1_2163(
      {stage51[111]},
      {stage51[116]}
   );
   gpc1_1 gpc1_1_2164(
      {stage51[112]},
      {stage51[117]}
   );
   gpc606_5 gpc606_5_2165(
      {stage53[112], stage53[113], stage53[114], stage53[115], stage53[116], stage53[117]},
      {stage55[107], stage55[108], stage55[109], stage55[110], stage55[111], stage55[112]},
      {stage57[114], stage56[146], stage55[114], stage54[126], stage53[120]}
   );
   gpc1_1 gpc1_1_2166(
      {stage54[115]},
      {stage54[127]}
   );
   gpc1_1 gpc1_1_2167(
      {stage54[116]},
      {stage54[128]}
   );
   gpc1_1 gpc1_1_2168(
      {stage54[117]},
      {stage54[129]}
   );
   gpc1_1 gpc1_1_2169(
      {stage54[118]},
      {stage54[130]}
   );
   gpc1_1 gpc1_1_2170(
      {stage54[119]},
      {stage54[131]}
   );
   gpc615_5 gpc615_5_2171(
      {stage54[120], stage54[121], stage54[122], stage54[123], stage54[124]},
      {stage55[113]},
      {stage56[130], stage56[131], stage56[132], stage56[133], stage56[134], stage56[135]},
      {stage58[121], stage57[115], stage56[147], stage55[115], stage54[132]}
   );
   gpc1_1 gpc1_1_2172(
      {stage56[136]},
      {stage56[148]}
   );
   gpc1_1 gpc1_1_2173(
      {stage56[137]},
      {stage56[149]}
   );
   gpc1_1 gpc1_1_2174(
      {stage56[138]},
      {stage56[150]}
   );
   gpc1_1 gpc1_1_2175(
      {stage56[139]},
      {stage56[151]}
   );
   gpc606_5 gpc606_5_2176(
      {stage56[140], stage56[141], stage56[142], stage56[143], stage56[144], stage56[145]},
      {stage58[114], stage58[115], stage58[116], stage58[117], stage58[118], stage58[119]},
      {stage60[131], stage59[130], stage58[122], stage57[116], stage56[152]}
   );
   gpc1_1 gpc1_1_2177(
      {stage57[108]},
      {stage57[117]}
   );
   gpc1_1 gpc1_1_2178(
      {stage57[109]},
      {stage57[118]}
   );
   gpc1_1 gpc1_1_2179(
      {stage57[110]},
      {stage57[119]}
   );
   gpc1_1 gpc1_1_2180(
      {stage57[111]},
      {stage57[120]}
   );
   gpc1_1 gpc1_1_2181(
      {stage57[112]},
      {stage57[121]}
   );
   gpc1_1 gpc1_1_2182(
      {stage57[113]},
      {stage57[122]}
   );
   gpc1_1 gpc1_1_2183(
      {stage58[120]},
      {stage58[123]}
   );
   gpc1_1 gpc1_1_2184(
      {stage59[121]},
      {stage59[131]}
   );
   gpc1_1 gpc1_1_2185(
      {stage59[122]},
      {stage59[132]}
   );
   gpc1_1 gpc1_1_2186(
      {stage59[123]},
      {stage59[133]}
   );
   gpc1_1 gpc1_1_2187(
      {stage59[124]},
      {stage59[134]}
   );
   gpc1_1 gpc1_1_2188(
      {stage59[125]},
      {stage59[135]}
   );
   gpc1_1 gpc1_1_2189(
      {stage59[126]},
      {stage59[136]}
   );
   gpc1_1 gpc1_1_2190(
      {stage59[127]},
      {stage59[137]}
   );
   gpc1_1 gpc1_1_2191(
      {stage59[128]},
      {stage59[138]}
   );
   gpc1_1 gpc1_1_2192(
      {stage59[129]},
      {stage59[139]}
   );
   gpc1_1 gpc1_1_2193(
      {stage60[117]},
      {stage60[132]}
   );
   gpc1_1 gpc1_1_2194(
      {stage60[118]},
      {stage60[133]}
   );
   gpc606_5 gpc606_5_2195(
      {stage60[119], stage60[120], stage60[121], stage60[122], stage60[123], stage60[124]},
      {stage62[110], stage62[111], stage62[112], stage62[113], stage62[114], stage62[115]},
      {stage64[43], stage63[115], stage62[128], stage61[133], stage60[134]}
   );
   gpc606_5 gpc606_5_2196(
      {stage60[125], stage60[126], stage60[127], stage60[128], stage60[129], stage60[130]},
      {stage62[116], stage62[117], stage62[118], stage62[119], stage62[120], stage62[121]},
      {stage64[44], stage63[116], stage62[129], stage61[134], stage60[135]}
   );
   gpc1_1 gpc1_1_2197(
      {stage61[125]},
      {stage61[135]}
   );
   gpc1_1 gpc1_1_2198(
      {stage61[126]},
      {stage61[136]}
   );
   gpc1_1 gpc1_1_2199(
      {stage61[127]},
      {stage61[137]}
   );
   gpc1_1 gpc1_1_2200(
      {stage61[128]},
      {stage61[138]}
   );
   gpc1_1 gpc1_1_2201(
      {stage61[129]},
      {stage61[139]}
   );
   gpc1_1 gpc1_1_2202(
      {stage61[130]},
      {stage61[140]}
   );
   gpc1_1 gpc1_1_2203(
      {stage61[131]},
      {stage61[141]}
   );
   gpc1_1 gpc1_1_2204(
      {stage61[132]},
      {stage61[142]}
   );
   gpc606_5 gpc606_5_2205(
      {stage62[122], stage62[123], stage62[124], stage62[125], stage62[126], stage62[127]},
      {stage64[31], stage64[32], stage64[33], stage64[34], stage64[35], stage64[36]},
      {stage66[7], stage65[27], stage64[45], stage63[117], stage62[130]}
   );
   gpc606_5 gpc606_5_2206(
      {stage63[110], stage63[111], stage63[112], stage63[113], stage63[114], 1'h0},
      {stage65[16], stage65[17], stage65[18], stage65[19], stage65[20], stage65[21]},
      {stage67[2], stage66[8], stage65[28], stage64[46], stage63[118]}
   );
   gpc1_1 gpc1_1_2207(
      {stage64[37]},
      {stage64[47]}
   );
   gpc135_4 gpc135_4_2208(
      {stage64[38], stage64[39], stage64[40], stage64[41], stage64[42]},
      {stage65[22], stage65[23], stage65[24]},
      {stage66[3]},
      {stage67[3], stage66[9], stage65[29], stage64[48]}
   );
   gpc1_1 gpc1_1_2209(
      {stage65[25]},
      {stage65[30]}
   );
   gpc1_1 gpc1_1_2210(
      {stage65[26]},
      {stage65[31]}
   );
   gpc1_1 gpc1_1_2211(
      {stage66[4]},
      {stage66[10]}
   );
   gpc1_1 gpc1_1_2212(
      {stage66[5]},
      {stage66[11]}
   );
   gpc1_1 gpc1_1_2213(
      {stage66[6]},
      {stage66[12]}
   );
   gpc1_1 gpc1_1_2214(
      {stage67[1]},
      {stage67[4]}
   );
   gpc1_1 gpc1_1_2215(
      {stage00[92]},
      {stage00[98]}
   );
   gpc2135_5 gpc2135_5_2216(
      {stage00[93], stage00[94], stage00[95], stage00[96], stage00[97]},
      {stage01[126], stage01[127], stage01[128]},
      {stage02[111]},
      {stage03[138], 1'h0},
      {stage04[124], stage03[139], stage02[117], stage01[129], stage00[99]}
   );
   gpc606_5 gpc606_5_2217(
      {stage02[112], stage02[113], stage02[114], stage02[115], stage02[116], 1'h0},
      {stage04[118], stage04[119], stage04[120], stage04[121], stage04[122], stage04[123]},
      {stage06[114], stage05[128], stage04[125], stage03[140], stage02[118]}
   );
   gpc606_5 gpc606_5_2218(
      {stage05[122], stage05[123], stage05[124], stage05[125], stage05[126], stage05[127]},
      {stage07[115], stage07[116], stage07[117], stage07[118], stage07[119], stage07[120]},
      {stage09[173], stage08[127], stage07[121], stage06[115], stage05[129]}
   );
   gpc1_1 gpc1_1_2219(
      {stage06[109]},
      {stage06[116]}
   );
   gpc1_1 gpc1_1_2220(
      {stage06[110]},
      {stage06[117]}
   );
   gpc1_1 gpc1_1_2221(
      {stage06[111]},
      {stage06[118]}
   );
   gpc1_1 gpc1_1_2222(
      {stage06[112]},
      {stage06[119]}
   );
   gpc1_1 gpc1_1_2223(
      {stage06[113]},
      {stage06[120]}
   );
   gpc615_5 gpc615_5_2224(
      {stage08[125], stage08[126], 1'h0, 1'h0, 1'h0},
      {stage09[167]},
      {stage10[139], stage10[140], stage10[141], stage10[142], stage10[143], stage10[144]},
      {stage12[151], stage11[158], stage10[145], stage09[174], stage08[128]}
   );
   gpc606_5 gpc606_5_2225(
      {stage09[168], stage09[169], stage09[170], stage09[171], stage09[172], 1'h0},
      {stage11[153], stage11[154], stage11[155], stage11[156], stage11[157], 1'h0},
      {stage13[138], stage12[152], stage11[159], stage10[146], stage09[175]}
   );
   gpc1_1 gpc1_1_2226(
      {stage12[143]},
      {stage12[153]}
   );
   gpc1_1 gpc1_1_2227(
      {stage12[144]},
      {stage12[154]}
   );
   gpc606_5 gpc606_5_2228(
      {stage12[145], stage12[146], stage12[147], stage12[148], stage12[149], stage12[150]},
      {stage14[110], stage14[111], stage14[112], stage14[113], stage14[114], stage14[115]},
      {stage16[113], stage15[166], stage14[116], stage13[139], stage12[155]}
   );
   gpc1406_5 gpc1406_5_2229(
      {stage13[126], stage13[127], stage13[128], stage13[129], stage13[130], stage13[131]},
      {stage15[156], stage15[157], stage15[158], stage15[159]},
      {stage16[111]},
      {stage17[153], stage16[114], stage15[167], stage14[117], stage13[140]}
   );
   gpc1406_5 gpc1406_5_2230(
      {stage13[132], stage13[133], stage13[134], stage13[135], stage13[136], stage13[137]},
      {stage15[160], stage15[161], stage15[162], stage15[163]},
      {stage16[112]},
      {stage17[154], stage16[115], stage15[168], stage14[118], stage13[141]}
   );
   gpc1_1 gpc1_1_2231(
      {stage15[164]},
      {stage15[169]}
   );
   gpc1_1 gpc1_1_2232(
      {stage15[165]},
      {stage15[170]}
   );
   gpc1_1 gpc1_1_2233(
      {stage17[149]},
      {stage17[155]}
   );
   gpc1_1 gpc1_1_2234(
      {stage17[150]},
      {stage17[156]}
   );
   gpc1_1 gpc1_1_2235(
      {stage17[151]},
      {stage17[157]}
   );
   gpc1_1 gpc1_1_2236(
      {stage17[152]},
      {stage17[158]}
   );
   gpc1_1 gpc1_1_2237(
      {stage18[120]},
      {stage18[127]}
   );
   gpc1_1 gpc1_1_2238(
      {stage18[121]},
      {stage18[128]}
   );
   gpc615_5 gpc615_5_2239(
      {stage18[122], stage18[123], stage18[124], stage18[125], stage18[126]},
      {stage19[122]},
      {stage20[147], stage20[148], stage20[149], stage20[150], stage20[151], stage20[152]},
      {stage22[120], stage21[118], stage20[154], stage19[131], stage18[129]}
   );
   gpc1_1 gpc1_1_2240(
      {stage19[123]},
      {stage19[132]}
   );
   gpc1_1 gpc1_1_2241(
      {stage19[124]},
      {stage19[133]}
   );
   gpc606_5 gpc606_5_2242(
      {stage19[125], stage19[126], stage19[127], stage19[128], stage19[129], stage19[130]},
      {stage21[112], stage21[113], stage21[114], stage21[115], stage21[116], stage21[117]},
      {stage23[141], stage22[121], stage21[119], stage20[155], stage19[134]}
   );
   gpc1_1 gpc1_1_2243(
      {stage20[153]},
      {stage20[156]}
   );
   gpc1_1 gpc1_1_2244(
      {stage22[113]},
      {stage22[122]}
   );
   gpc1_1 gpc1_1_2245(
      {stage22[114]},
      {stage22[123]}
   );
   gpc615_5 gpc615_5_2246(
      {stage22[115], stage22[116], stage22[117], stage22[118], stage22[119]},
      {stage23[135]},
      {stage24[117], stage24[118], stage24[119], stage24[120], stage24[121], stage24[122]},
      {stage26[112], stage25[137], stage24[124], stage23[142], stage22[124]}
   );
   gpc1_1 gpc1_1_2247(
      {stage23[136]},
      {stage23[143]}
   );
   gpc1_1 gpc1_1_2248(
      {stage23[137]},
      {stage23[144]}
   );
   gpc1_1 gpc1_1_2249(
      {stage23[138]},
      {stage23[145]}
   );
   gpc1_1 gpc1_1_2250(
      {stage23[139]},
      {stage23[146]}
   );
   gpc1_1 gpc1_1_2251(
      {stage23[140]},
      {stage23[147]}
   );
   gpc1_1 gpc1_1_2252(
      {stage24[123]},
      {stage24[125]}
   );
   gpc606_5 gpc606_5_2253(
      {stage25[132], stage25[133], stage25[134], stage25[135], stage25[136], 1'h0},
      {stage27[136], stage27[137], stage27[138], stage27[139], stage27[140], stage27[141]},
      {stage29[114], stage28[145], stage27[147], stage26[113], stage25[138]}
   );
   gpc1_1 gpc1_1_2254(
      {stage26[103]},
      {stage26[114]}
   );
   gpc1_1 gpc1_1_2255(
      {stage26[104]},
      {stage26[115]}
   );
   gpc7_3 gpc7_3_2256(
      {stage26[105], stage26[106], stage26[107], stage26[108], stage26[109], stage26[110], stage26[111]},
      {stage28[146], stage27[148], stage26[116]}
   );
   gpc615_5 gpc615_5_2257(
      {stage27[142], stage27[143], stage27[144], stage27[145], stage27[146]},
      {stage28[138]},
      {stage29[107], stage29[108], stage29[109], stage29[110], stage29[111], stage29[112]},
      {stage31[126], stage30[135], stage29[115], stage28[147], stage27[149]}
   );
   gpc1_1 gpc1_1_2258(
      {stage28[139]},
      {stage28[148]}
   );
   gpc615_5 gpc615_5_2259(
      {stage28[140], stage28[141], stage28[142], stage28[143], stage28[144]},
      {stage29[113]},
      {stage30[129], stage30[130], stage30[131], stage30[132], stage30[133], stage30[134]},
      {stage32[114], stage31[127], stage30[136], stage29[116], stage28[149]}
   );
   gpc135_4 gpc135_4_2260(
      {stage31[122], stage31[123], stage31[124], stage31[125], 1'h0},
      {stage32[111], stage32[112], stage32[113]},
      {stage33[110]},
      {stage34[117], stage33[113], stage32[115], stage31[128]}
   );
   gpc1343_5 gpc1343_5_2261(
      {stage33[111], stage33[112], 1'h0},
      {stage34[109], stage34[110], stage34[111], stage34[112]},
      {stage35[112], stage35[113], stage35[114]},
      {stage36[132]},
      {stage37[126], stage36[143], stage35[115], stage34[118], stage33[114]}
   );
   gpc1_1 gpc1_1_2262(
      {stage34[113]},
      {stage34[119]}
   );
   gpc1_1 gpc1_1_2263(
      {stage34[114]},
      {stage34[120]}
   );
   gpc1_1 gpc1_1_2264(
      {stage34[115]},
      {stage34[121]}
   );
   gpc1_1 gpc1_1_2265(
      {stage34[116]},
      {stage34[122]}
   );
   gpc1_1 gpc1_1_2266(
      {stage36[133]},
      {stage36[144]}
   );
   gpc1_1 gpc1_1_2267(
      {stage36[134]},
      {stage36[145]}
   );
   gpc1_1 gpc1_1_2268(
      {stage36[135]},
      {stage36[146]}
   );
   gpc1_1 gpc1_1_2269(
      {stage36[136]},
      {stage36[147]}
   );
   gpc606_5 gpc606_5_2270(
      {stage36[137], stage36[138], stage36[139], stage36[140], stage36[141], stage36[142]},
      {stage38[114], stage38[115], stage38[116], stage38[117], stage38[118], 1'h0},
      {stage40[137], stage39[116], stage38[119], stage37[127], stage36[148]}
   );
   gpc606_5 gpc606_5_2271(
      {stage37[120], stage37[121], stage37[122], stage37[123], stage37[124], stage37[125]},
      {stage39[109], stage39[110], stage39[111], stage39[112], stage39[113], stage39[114]},
      {stage41[144], stage40[138], stage39[117], stage38[120], stage37[128]}
   );
   gpc1_1 gpc1_1_2272(
      {stage39[115]},
      {stage39[118]}
   );
   gpc1_1 gpc1_1_2273(
      {stage40[131]},
      {stage40[139]}
   );
   gpc1_1 gpc1_1_2274(
      {stage40[132]},
      {stage40[140]}
   );
   gpc1_1 gpc1_1_2275(
      {stage40[133]},
      {stage40[141]}
   );
   gpc1343_5 gpc1343_5_2276(
      {stage40[134], stage40[135], stage40[136]},
      {stage41[139], stage41[140], stage41[141], stage41[142]},
      {stage42[137], stage42[138], stage42[139]},
      {stage43[151]},
      {stage44[122], stage43[157], stage42[141], stage41[145], stage40[142]}
   );
   gpc1_1 gpc1_1_2277(
      {stage41[143]},
      {stage41[146]}
   );
   gpc1_1 gpc1_1_2278(
      {stage42[140]},
      {stage42[142]}
   );
   gpc615_5 gpc615_5_2279(
      {stage43[152], stage43[153], stage43[154], stage43[155], stage43[156]},
      {stage44[117]},
      {stage45[135], stage45[136], stage45[137], stage45[138], stage45[139], stage45[140]},
      {stage47[134], stage46[130], stage45[141], stage44[123], stage43[158]}
   );
   gpc1_1 gpc1_1_2280(
      {stage44[118]},
      {stage44[124]}
   );
   gpc1_1 gpc1_1_2281(
      {stage44[119]},
      {stage44[125]}
   );
   gpc1_1 gpc1_1_2282(
      {stage44[120]},
      {stage44[126]}
   );
   gpc1_1 gpc1_1_2283(
      {stage44[121]},
      {stage44[127]}
   );
   gpc1_1 gpc1_1_2284(
      {stage46[125]},
      {stage46[131]}
   );
   gpc1_1 gpc1_1_2285(
      {stage46[126]},
      {stage46[132]}
   );
   gpc1_1 gpc1_1_2286(
      {stage46[127]},
      {stage46[133]}
   );
   gpc1_1 gpc1_1_2287(
      {stage46[128]},
      {stage46[134]}
   );
   gpc1_1 gpc1_1_2288(
      {stage46[129]},
      {stage46[135]}
   );
   gpc135_4 gpc135_4_2289(
      {stage47[126], stage47[127], stage47[128], stage47[129], stage47[130]},
      {stage48[124], stage48[125], stage48[126]},
      {stage49[133]},
      {stage50[121], stage49[145], stage48[128], stage47[135]}
   );
   gpc135_4 gpc135_4_2290(
      {stage47[131], stage47[132], stage47[133], 1'h0, 1'h0},
      {stage48[127], 1'h0, 1'h0},
      {stage49[134]},
      {stage50[122], stage49[146], stage48[129], stage47[136]}
   );
   gpc1_1 gpc1_1_2291(
      {stage49[135]},
      {stage49[147]}
   );
   gpc1_1 gpc1_1_2292(
      {stage49[136]},
      {stage49[148]}
   );
   gpc1_1 gpc1_1_2293(
      {stage49[137]},
      {stage49[149]}
   );
   gpc1_1 gpc1_1_2294(
      {stage49[138]},
      {stage49[150]}
   );
   gpc606_5 gpc606_5_2295(
      {stage49[139], stage49[140], stage49[141], stage49[142], stage49[143], stage49[144]},
      {stage51[113], stage51[114], stage51[115], stage51[116], stage51[117], 1'h0},
      {stage53[121], stage52[118], stage51[118], stage50[123], stage49[151]}
   );
   gpc7_3 gpc7_3_2296(
      {stage50[116], stage50[117], stage50[118], stage50[119], stage50[120], 1'h0, 1'h0},
      {stage52[119], stage51[119], stage50[124]}
   );
   gpc1_1 gpc1_1_2297(
      {stage52[116]},
      {stage52[120]}
   );
   gpc1_1 gpc1_1_2298(
      {stage52[117]},
      {stage52[121]}
   );
   gpc1_1 gpc1_1_2299(
      {stage53[118]},
      {stage53[122]}
   );
   gpc1_1 gpc1_1_2300(
      {stage53[119]},
      {stage53[123]}
   );
   gpc1_1 gpc1_1_2301(
      {stage53[120]},
      {stage53[124]}
   );
   gpc1_1 gpc1_1_2302(
      {stage54[125]},
      {stage54[133]}
   );
   gpc1_1 gpc1_1_2303(
      {stage54[126]},
      {stage54[134]}
   );
   gpc1_1 gpc1_1_2304(
      {stage54[127]},
      {stage54[135]}
   );
   gpc1_1 gpc1_1_2305(
      {stage54[128]},
      {stage54[136]}
   );
   gpc1_1 gpc1_1_2306(
      {stage54[129]},
      {stage54[137]}
   );
   gpc623_5 gpc623_5_2307(
      {stage54[130], stage54[131], stage54[132]},
      {stage55[114], stage55[115]},
      {stage56[146], stage56[147], stage56[148], stage56[149], stage56[150], stage56[151]},
      {stage58[124], stage57[123], stage56[153], stage55[116], stage54[138]}
   );
   gpc1_1 gpc1_1_2308(
      {stage56[152]},
      {stage56[154]}
   );
   gpc1_1 gpc1_1_2309(
      {stage57[114]},
      {stage57[124]}
   );
   gpc1_1 gpc1_1_2310(
      {stage57[115]},
      {stage57[125]}
   );
   gpc1_1 gpc1_1_2311(
      {stage57[116]},
      {stage57[126]}
   );
   gpc606_5 gpc606_5_2312(
      {stage57[117], stage57[118], stage57[119], stage57[120], stage57[121], stage57[122]},
      {stage59[130], stage59[131], stage59[132], stage59[133], stage59[134], stage59[135]},
      {stage61[143], stage60[136], stage59[140], stage58[125], stage57[127]}
   );
   gpc623_5 gpc623_5_2313(
      {stage58[121], stage58[122], stage58[123]},
      {stage59[136], stage59[137]},
      {stage60[131], stage60[132], stage60[133], stage60[134], stage60[135], 1'h0},
      {stage62[131], stage61[144], stage60[137], stage59[141], stage58[126]}
   );
   gpc1_1 gpc1_1_2314(
      {stage59[138]},
      {stage59[142]}
   );
   gpc1_1 gpc1_1_2315(
      {stage59[139]},
      {stage59[143]}
   );
   gpc1_1 gpc1_1_2316(
      {stage61[133]},
      {stage61[145]}
   );
   gpc1_1 gpc1_1_2317(
      {stage61[134]},
      {stage61[146]}
   );
   gpc1_1 gpc1_1_2318(
      {stage61[135]},
      {stage61[147]}
   );
   gpc1_1 gpc1_1_2319(
      {stage61[136]},
      {stage61[148]}
   );
   gpc606_5 gpc606_5_2320(
      {stage61[137], stage61[138], stage61[139], stage61[140], stage61[141], stage61[142]},
      {stage63[115], stage63[116], stage63[117], stage63[118], 1'h0, 1'h0},
      {stage65[32], stage64[49], stage63[119], stage62[132], stage61[149]}
   );
   gpc1_1 gpc1_1_2321(
      {stage62[128]},
      {stage62[133]}
   );
   gpc1_1 gpc1_1_2322(
      {stage62[129]},
      {stage62[134]}
   );
   gpc1_1 gpc1_1_2323(
      {stage62[130]},
      {stage62[135]}
   );
   gpc1406_5 gpc1406_5_2324(
      {stage64[43], stage64[44], stage64[45], stage64[46], stage64[47], stage64[48]},
      {stage66[7], stage66[8], stage66[9], stage66[10]},
      {stage67[2]},
      {stage68[0], stage67[5], stage66[13], stage65[33], stage64[50]}
   );
   gpc1_1 gpc1_1_2325(
      {stage65[27]},
      {stage65[34]}
   );
   gpc1_1 gpc1_1_2326(
      {stage65[28]},
      {stage65[35]}
   );
   gpc1343_5 gpc1343_5_2327(
      {stage65[29], stage65[30], stage65[31]},
      {stage66[11], stage66[12], 1'h0, 1'h0},
      {stage67[3], stage67[4], 1'h0},
      {1'h0},
      {stage69[0], stage68[1], stage67[6], stage66[14], stage65[36]}
   );
   gpc1_1 gpc1_1_2328(
      {stage00[98]},
      {stage00[100]}
   );
   gpc1_1 gpc1_1_2329(
      {stage00[99]},
      {stage00[101]}
   );
   gpc1_1 gpc1_1_2330(
      {stage01[129]},
      {stage01[130]}
   );
   gpc1_1 gpc1_1_2331(
      {stage02[117]},
      {stage02[119]}
   );
   gpc1_1 gpc1_1_2332(
      {stage02[118]},
      {stage02[120]}
   );
   gpc1_1 gpc1_1_2333(
      {stage03[139]},
      {stage03[141]}
   );
   gpc1_1 gpc1_1_2334(
      {stage03[140]},
      {stage03[142]}
   );
   gpc1_1 gpc1_1_2335(
      {stage04[124]},
      {stage04[126]}
   );
   gpc1_1 gpc1_1_2336(
      {stage04[125]},
      {stage04[127]}
   );
   gpc1_1 gpc1_1_2337(
      {stage05[128]},
      {stage05[130]}
   );
   gpc1_1 gpc1_1_2338(
      {stage05[129]},
      {stage05[131]}
   );
   gpc1_1 gpc1_1_2339(
      {stage06[114]},
      {stage06[121]}
   );
   gpc606_5 gpc606_5_2340(
      {stage06[115], stage06[116], stage06[117], stage06[118], stage06[119], stage06[120]},
      {stage08[127], stage08[128], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage10[147], stage09[176], stage08[129], stage07[122], stage06[122]}
   );
   gpc1_1 gpc1_1_2341(
      {stage07[121]},
      {stage07[123]}
   );
   gpc135_4 gpc135_4_2342(
      {stage09[173], stage09[174], stage09[175], 1'h0, 1'h0},
      {stage10[145], stage10[146], 1'h0},
      {stage11[158]},
      {stage12[156], stage11[160], stage10[148], stage09[177]}
   );
   gpc1_1 gpc1_1_2343(
      {stage11[159]},
      {stage11[161]}
   );
   gpc7_3 gpc7_3_2344(
      {stage12[151], stage12[152], stage12[153], stage12[154], stage12[155], 1'h0, 1'h0},
      {stage14[119], stage13[142], stage12[157]}
   );
   gpc2135_5 gpc2135_5_2345(
      {stage13[138], stage13[139], stage13[140], stage13[141], 1'h0},
      {stage14[116], stage14[117], stage14[118]},
      {stage15[166]},
      {stage16[113], stage16[114]},
      {stage17[159], stage16[116], stage15[171], stage14[120], stage13[143]}
   );
   gpc615_5 gpc615_5_2346(
      {stage15[167], stage15[168], stage15[169], stage15[170], 1'h0},
      {stage16[115]},
      {stage17[153], stage17[154], stage17[155], stage17[156], stage17[157], stage17[158]},
      {stage19[135], stage18[130], stage17[160], stage16[117], stage15[172]}
   );
   gpc1343_5 gpc1343_5_2347(
      {stage18[127], stage18[128], stage18[129]},
      {stage19[131], stage19[132], stage19[133], stage19[134]},
      {stage20[154], stage20[155], stage20[156]},
      {stage21[118]},
      {stage22[125], stage21[120], stage20[157], stage19[136], stage18[131]}
   );
   gpc1_1 gpc1_1_2348(
      {stage21[119]},
      {stage21[121]}
   );
   gpc215_4 gpc215_4_2349(
      {stage22[120], stage22[121], stage22[122], stage22[123], stage22[124]},
      {stage23[141]},
      {stage24[124], stage24[125]},
      {stage25[139], stage24[126], stage23[148], stage22[126]}
   );
   gpc207_4 gpc207_4_2350(
      {stage23[142], stage23[143], stage23[144], stage23[145], stage23[146], stage23[147], 1'h0},
      {stage25[137], stage25[138]},
      {stage26[117], stage25[140], stage24[127], stage23[149]}
   );
   gpc615_5 gpc615_5_2351(
      {stage26[112], stage26[113], stage26[114], stage26[115], stage26[116]},
      {stage27[147]},
      {stage28[145], stage28[146], stage28[147], stage28[148], stage28[149], 1'h0},
      {stage30[137], stage29[117], stage28[150], stage27[150], stage26[118]}
   );
   gpc3_2 gpc3_2_2352(
      {stage27[148], stage27[149], 1'h0},
      {stage28[151], stage27[151]}
   );
   gpc1343_5 gpc1343_5_2353(
      {stage29[114], stage29[115], stage29[116]},
      {stage30[135], stage30[136], 1'h0, 1'h0},
      {stage31[126], stage31[127], stage31[128]},
      {stage32[114]},
      {stage33[115], stage32[116], stage31[129], stage30[138], stage29[118]}
   );
   gpc623_5 gpc623_5_2354(
      {stage32[115], 1'h0, 1'h0},
      {stage33[113], stage33[114]},
      {stage34[117], stage34[118], stage34[119], stage34[120], stage34[121], stage34[122]},
      {stage36[149], stage35[116], stage34[123], stage33[116], stage32[117]}
   );
   gpc1_1 gpc1_1_2355(
      {stage35[115]},
      {stage35[117]}
   );
   gpc207_4 gpc207_4_2356(
      {stage36[143], stage36[144], stage36[145], stage36[146], stage36[147], stage36[148], 1'h0},
      {stage38[119], stage38[120]},
      {stage39[119], stage38[121], stage37[129], stage36[150]}
   );
   gpc3_2 gpc3_2_2357(
      {stage37[126], stage37[127], stage37[128]},
      {stage38[122], stage37[130]}
   );
   gpc3_2 gpc3_2_2358(
      {stage39[116], stage39[117], stage39[118]},
      {stage40[143], stage39[120]}
   );
   gpc7_3 gpc7_3_2359(
      {stage40[137], stage40[138], stage40[139], stage40[140], stage40[141], stage40[142], 1'h0},
      {stage42[143], stage41[147], stage40[144]}
   );
   gpc135_4 gpc135_4_2360(
      {stage41[144], stage41[145], stage41[146], 1'h0, 1'h0},
      {stage42[141], stage42[142], 1'h0},
      {stage43[157]},
      {stage44[128], stage43[159], stage42[144], stage41[148]}
   );
   gpc1_1 gpc1_1_2361(
      {stage43[158]},
      {stage43[160]}
   );
   gpc606_5 gpc606_5_2362(
      {stage44[122], stage44[123], stage44[124], stage44[125], stage44[126], stage44[127]},
      {stage46[130], stage46[131], stage46[132], stage46[133], stage46[134], stage46[135]},
      {stage48[130], stage47[137], stage46[136], stage45[142], stage44[129]}
   );
   gpc1_1 gpc1_1_2363(
      {stage45[141]},
      {stage45[143]}
   );
   gpc623_5 gpc623_5_2364(
      {stage47[134], stage47[135], stage47[136]},
      {stage48[128], stage48[129]},
      {stage49[145], stage49[146], stage49[147], stage49[148], stage49[149], stage49[150]},
      {stage51[120], stage50[125], stage49[152], stage48[131], stage47[138]}
   );
   gpc1_1 gpc1_1_2365(
      {stage49[151]},
      {stage49[153]}
   );
   gpc2135_5 gpc2135_5_2366(
      {stage50[121], stage50[122], stage50[123], stage50[124], 1'h0},
      {stage51[118], stage51[119], 1'h0},
      {stage52[118]},
      {stage53[121], stage53[122]},
      {stage54[139], stage53[125], stage52[122], stage51[121], stage50[126]}
   );
   gpc623_5 gpc623_5_2367(
      {stage52[119], stage52[120], stage52[121]},
      {stage53[123], stage53[124]},
      {stage54[133], stage54[134], stage54[135], stage54[136], stage54[137], stage54[138]},
      {stage56[155], stage55[117], stage54[140], stage53[126], stage52[123]}
   );
   gpc1_1 gpc1_1_2368(
      {stage55[116]},
      {stage55[118]}
   );
   gpc1343_5 gpc1343_5_2369(
      {stage56[153], stage56[154], 1'h0},
      {stage57[123], stage57[124], stage57[125], stage57[126]},
      {stage58[124], stage58[125], stage58[126]},
      {stage59[140]},
      {stage60[138], stage59[144], stage58[127], stage57[128], stage56[156]}
   );
   gpc1_1 gpc1_1_2370(
      {stage57[127]},
      {stage57[129]}
   );
   gpc623_5 gpc623_5_2371(
      {stage59[141], stage59[142], stage59[143]},
      {stage60[136], stage60[137]},
      {stage61[143], stage61[144], stage61[145], stage61[146], stage61[147], stage61[148]},
      {stage63[120], stage62[136], stage61[150], stage60[139], stage59[145]}
   );
   gpc1_1 gpc1_1_2372(
      {stage61[149]},
      {stage61[151]}
   );
   gpc215_4 gpc215_4_2373(
      {stage62[131], stage62[132], stage62[133], stage62[134], stage62[135]},
      {stage63[119]},
      {stage64[49], stage64[50]},
      {stage65[37], stage64[51], stage63[121], stage62[137]}
   );
   gpc207_4 gpc207_4_2374(
      {stage65[32], stage65[33], stage65[34], stage65[35], stage65[36], 1'h0, 1'h0},
      {stage67[5], stage67[6]},
      {stage68[2], stage67[7], stage66[15], stage65[38]}
   );
   gpc606_5 gpc606_5_2375(
      {stage66[13], stage66[14], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage68[0], stage68[1], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage70[0], stage69[1], stage68[3], stage67[8], stage66[16]}
   );
   gpc1_1 gpc1_1_2376(
      {stage69[0]},
      {stage69[2]}
   );
endmodule

module behavioral_tester();
   reg [63:0] src00;
   reg [63:0] src01;
   reg [63:0] src02;
   reg [63:0] src03;
   reg [63:0] src04;
   reg [63:0] src05;
   reg [63:0] src06;
   reg [63:0] src07;
   reg [63:0] src08;
   reg [63:0] src09;
   reg [63:0] src10;
   reg [63:0] src11;
   reg [63:0] src12;
   reg [63:0] src13;
   reg [63:0] src14;
   reg [63:0] src15;
   reg [63:0] src16;
   reg [63:0] src17;
   reg [63:0] src18;
   reg [63:0] src19;
   reg [63:0] src20;
   reg [63:0] src21;
   reg [63:0] src22;
   reg [63:0] src23;
   reg [63:0] src24;
   reg [63:0] src25;
   reg [63:0] src26;
   reg [63:0] src27;
   reg [63:0] src28;
   reg [63:0] src29;
   reg [63:0] src30;
   reg [63:0] src31;
   reg [63:0] src32;
   reg [63:0] src33;
   reg [63:0] src34;
   reg [63:0] src35;
   reg [63:0] src36;
   reg [63:0] src37;
   reg [63:0] src38;
   reg [63:0] src39;
   reg [63:0] src40;
   reg [63:0] src41;
   reg [63:0] src42;
   reg [63:0] src43;
   reg [63:0] src44;
   reg [63:0] src45;
   reg [63:0] src46;
   reg [63:0] src47;
   reg [63:0] src48;
   reg [63:0] src49;
   reg [63:0] src50;
   reg [63:0] src51;
   reg [63:0] src52;
   reg [63:0] src53;
   reg [63:0] src54;
   reg [63:0] src55;
   reg [63:0] src56;
   reg [63:0] src57;
   reg [63:0] src58;
   reg [63:0] src59;
   reg [63:0] src60;
   reg [63:0] src61;
   reg [63:0] src62;
   reg [63:0] src63;
   wire [1:0] dst00;
   wire [0:0] dst01;
   wire [1:0] dst02;
   wire [1:0] dst03;
   wire [1:0] dst04;
   wire [1:0] dst05;
   wire [1:0] dst06;
   wire [1:0] dst07;
   wire [0:0] dst08;
   wire [1:0] dst09;
   wire [1:0] dst10;
   wire [1:0] dst11;
   wire [1:0] dst12;
   wire [1:0] dst13;
   wire [1:0] dst14;
   wire [1:0] dst15;
   wire [1:0] dst16;
   wire [1:0] dst17;
   wire [1:0] dst18;
   wire [1:0] dst19;
   wire [0:0] dst20;
   wire [1:0] dst21;
   wire [1:0] dst22;
   wire [1:0] dst23;
   wire [1:0] dst24;
   wire [1:0] dst25;
   wire [1:0] dst26;
   wire [1:0] dst27;
   wire [1:0] dst28;
   wire [1:0] dst29;
   wire [1:0] dst30;
   wire [0:0] dst31;
   wire [1:0] dst32;
   wire [1:0] dst33;
   wire [0:0] dst34;
   wire [1:0] dst35;
   wire [1:0] dst36;
   wire [1:0] dst37;
   wire [1:0] dst38;
   wire [1:0] dst39;
   wire [1:0] dst40;
   wire [1:0] dst41;
   wire [1:0] dst42;
   wire [1:0] dst43;
   wire [1:0] dst44;
   wire [1:0] dst45;
   wire [0:0] dst46;
   wire [1:0] dst47;
   wire [1:0] dst48;
   wire [1:0] dst49;
   wire [1:0] dst50;
   wire [1:0] dst51;
   wire [1:0] dst52;
   wire [1:0] dst53;
   wire [1:0] dst54;
   wire [1:0] dst55;
   wire [1:0] dst56;
   wire [1:0] dst57;
   wire [0:0] dst58;
   wire [1:0] dst59;
   wire [1:0] dst60;
   wire [1:0] dst61;
   wire [1:0] dst62;
   wire [1:0] dst63;
   wire [0:0] dst64;
   wire [1:0] dst65;
   wire [1:0] dst66;
   wire [1:0] dst67;
   wire [1:0] dst68;
   wire [1:0] dst69;
   wire [0:0] dst70;
   wire [71:0] srcsum;
   wire [71:0] dstsum;
   wire test;
   assign srcsum =
      (src00[0] << 0) +
      (src00[1] << 0) +
      (src00[2] << 0) +
      (src00[3] << 0) +
      (src00[4] << 0) +
      (src00[5] << 0) +
      (src00[6] << 0) +
      (src00[7] << 0) +
      (src00[8] << 0) +
      (src00[9] << 0) +
      (src00[10] << 0) +
      (src00[11] << 0) +
      (src00[12] << 0) +
      (src00[13] << 0) +
      (src00[14] << 0) +
      (src00[15] << 0) +
      (src00[16] << 0) +
      (src00[17] << 0) +
      (src00[18] << 0) +
      (src00[19] << 0) +
      (src00[20] << 0) +
      (src00[21] << 0) +
      (src00[22] << 0) +
      (src00[23] << 0) +
      (src00[24] << 0) +
      (src00[25] << 0) +
      (src00[26] << 0) +
      (src00[27] << 0) +
      (src00[28] << 0) +
      (src00[29] << 0) +
      (src00[30] << 0) +
      (src00[31] << 0) +
      (src00[32] << 0) +
      (src00[33] << 0) +
      (src00[34] << 0) +
      (src00[35] << 0) +
      (src00[36] << 0) +
      (src00[37] << 0) +
      (src00[38] << 0) +
      (src00[39] << 0) +
      (src00[40] << 0) +
      (src00[41] << 0) +
      (src00[42] << 0) +
      (src00[43] << 0) +
      (src00[44] << 0) +
      (src00[45] << 0) +
      (src00[46] << 0) +
      (src00[47] << 0) +
      (src00[48] << 0) +
      (src00[49] << 0) +
      (src00[50] << 0) +
      (src00[51] << 0) +
      (src00[52] << 0) +
      (src00[53] << 0) +
      (src00[54] << 0) +
      (src00[55] << 0) +
      (src00[56] << 0) +
      (src00[57] << 0) +
      (src00[58] << 0) +
      (src00[59] << 0) +
      (src00[60] << 0) +
      (src00[61] << 0) +
      (src00[62] << 0) +
      (src00[63] << 0) +
      (src01[0] << 1) +
      (src01[1] << 1) +
      (src01[2] << 1) +
      (src01[3] << 1) +
      (src01[4] << 1) +
      (src01[5] << 1) +
      (src01[6] << 1) +
      (src01[7] << 1) +
      (src01[8] << 1) +
      (src01[9] << 1) +
      (src01[10] << 1) +
      (src01[11] << 1) +
      (src01[12] << 1) +
      (src01[13] << 1) +
      (src01[14] << 1) +
      (src01[15] << 1) +
      (src01[16] << 1) +
      (src01[17] << 1) +
      (src01[18] << 1) +
      (src01[19] << 1) +
      (src01[20] << 1) +
      (src01[21] << 1) +
      (src01[22] << 1) +
      (src01[23] << 1) +
      (src01[24] << 1) +
      (src01[25] << 1) +
      (src01[26] << 1) +
      (src01[27] << 1) +
      (src01[28] << 1) +
      (src01[29] << 1) +
      (src01[30] << 1) +
      (src01[31] << 1) +
      (src01[32] << 1) +
      (src01[33] << 1) +
      (src01[34] << 1) +
      (src01[35] << 1) +
      (src01[36] << 1) +
      (src01[37] << 1) +
      (src01[38] << 1) +
      (src01[39] << 1) +
      (src01[40] << 1) +
      (src01[41] << 1) +
      (src01[42] << 1) +
      (src01[43] << 1) +
      (src01[44] << 1) +
      (src01[45] << 1) +
      (src01[46] << 1) +
      (src01[47] << 1) +
      (src01[48] << 1) +
      (src01[49] << 1) +
      (src01[50] << 1) +
      (src01[51] << 1) +
      (src01[52] << 1) +
      (src01[53] << 1) +
      (src01[54] << 1) +
      (src01[55] << 1) +
      (src01[56] << 1) +
      (src01[57] << 1) +
      (src01[58] << 1) +
      (src01[59] << 1) +
      (src01[60] << 1) +
      (src01[61] << 1) +
      (src01[62] << 1) +
      (src01[63] << 1) +
      (src02[0] << 2) +
      (src02[1] << 2) +
      (src02[2] << 2) +
      (src02[3] << 2) +
      (src02[4] << 2) +
      (src02[5] << 2) +
      (src02[6] << 2) +
      (src02[7] << 2) +
      (src02[8] << 2) +
      (src02[9] << 2) +
      (src02[10] << 2) +
      (src02[11] << 2) +
      (src02[12] << 2) +
      (src02[13] << 2) +
      (src02[14] << 2) +
      (src02[15] << 2) +
      (src02[16] << 2) +
      (src02[17] << 2) +
      (src02[18] << 2) +
      (src02[19] << 2) +
      (src02[20] << 2) +
      (src02[21] << 2) +
      (src02[22] << 2) +
      (src02[23] << 2) +
      (src02[24] << 2) +
      (src02[25] << 2) +
      (src02[26] << 2) +
      (src02[27] << 2) +
      (src02[28] << 2) +
      (src02[29] << 2) +
      (src02[30] << 2) +
      (src02[31] << 2) +
      (src02[32] << 2) +
      (src02[33] << 2) +
      (src02[34] << 2) +
      (src02[35] << 2) +
      (src02[36] << 2) +
      (src02[37] << 2) +
      (src02[38] << 2) +
      (src02[39] << 2) +
      (src02[40] << 2) +
      (src02[41] << 2) +
      (src02[42] << 2) +
      (src02[43] << 2) +
      (src02[44] << 2) +
      (src02[45] << 2) +
      (src02[46] << 2) +
      (src02[47] << 2) +
      (src02[48] << 2) +
      (src02[49] << 2) +
      (src02[50] << 2) +
      (src02[51] << 2) +
      (src02[52] << 2) +
      (src02[53] << 2) +
      (src02[54] << 2) +
      (src02[55] << 2) +
      (src02[56] << 2) +
      (src02[57] << 2) +
      (src02[58] << 2) +
      (src02[59] << 2) +
      (src02[60] << 2) +
      (src02[61] << 2) +
      (src02[62] << 2) +
      (src02[63] << 2) +
      (src03[0] << 3) +
      (src03[1] << 3) +
      (src03[2] << 3) +
      (src03[3] << 3) +
      (src03[4] << 3) +
      (src03[5] << 3) +
      (src03[6] << 3) +
      (src03[7] << 3) +
      (src03[8] << 3) +
      (src03[9] << 3) +
      (src03[10] << 3) +
      (src03[11] << 3) +
      (src03[12] << 3) +
      (src03[13] << 3) +
      (src03[14] << 3) +
      (src03[15] << 3) +
      (src03[16] << 3) +
      (src03[17] << 3) +
      (src03[18] << 3) +
      (src03[19] << 3) +
      (src03[20] << 3) +
      (src03[21] << 3) +
      (src03[22] << 3) +
      (src03[23] << 3) +
      (src03[24] << 3) +
      (src03[25] << 3) +
      (src03[26] << 3) +
      (src03[27] << 3) +
      (src03[28] << 3) +
      (src03[29] << 3) +
      (src03[30] << 3) +
      (src03[31] << 3) +
      (src03[32] << 3) +
      (src03[33] << 3) +
      (src03[34] << 3) +
      (src03[35] << 3) +
      (src03[36] << 3) +
      (src03[37] << 3) +
      (src03[38] << 3) +
      (src03[39] << 3) +
      (src03[40] << 3) +
      (src03[41] << 3) +
      (src03[42] << 3) +
      (src03[43] << 3) +
      (src03[44] << 3) +
      (src03[45] << 3) +
      (src03[46] << 3) +
      (src03[47] << 3) +
      (src03[48] << 3) +
      (src03[49] << 3) +
      (src03[50] << 3) +
      (src03[51] << 3) +
      (src03[52] << 3) +
      (src03[53] << 3) +
      (src03[54] << 3) +
      (src03[55] << 3) +
      (src03[56] << 3) +
      (src03[57] << 3) +
      (src03[58] << 3) +
      (src03[59] << 3) +
      (src03[60] << 3) +
      (src03[61] << 3) +
      (src03[62] << 3) +
      (src03[63] << 3) +
      (src04[0] << 4) +
      (src04[1] << 4) +
      (src04[2] << 4) +
      (src04[3] << 4) +
      (src04[4] << 4) +
      (src04[5] << 4) +
      (src04[6] << 4) +
      (src04[7] << 4) +
      (src04[8] << 4) +
      (src04[9] << 4) +
      (src04[10] << 4) +
      (src04[11] << 4) +
      (src04[12] << 4) +
      (src04[13] << 4) +
      (src04[14] << 4) +
      (src04[15] << 4) +
      (src04[16] << 4) +
      (src04[17] << 4) +
      (src04[18] << 4) +
      (src04[19] << 4) +
      (src04[20] << 4) +
      (src04[21] << 4) +
      (src04[22] << 4) +
      (src04[23] << 4) +
      (src04[24] << 4) +
      (src04[25] << 4) +
      (src04[26] << 4) +
      (src04[27] << 4) +
      (src04[28] << 4) +
      (src04[29] << 4) +
      (src04[30] << 4) +
      (src04[31] << 4) +
      (src04[32] << 4) +
      (src04[33] << 4) +
      (src04[34] << 4) +
      (src04[35] << 4) +
      (src04[36] << 4) +
      (src04[37] << 4) +
      (src04[38] << 4) +
      (src04[39] << 4) +
      (src04[40] << 4) +
      (src04[41] << 4) +
      (src04[42] << 4) +
      (src04[43] << 4) +
      (src04[44] << 4) +
      (src04[45] << 4) +
      (src04[46] << 4) +
      (src04[47] << 4) +
      (src04[48] << 4) +
      (src04[49] << 4) +
      (src04[50] << 4) +
      (src04[51] << 4) +
      (src04[52] << 4) +
      (src04[53] << 4) +
      (src04[54] << 4) +
      (src04[55] << 4) +
      (src04[56] << 4) +
      (src04[57] << 4) +
      (src04[58] << 4) +
      (src04[59] << 4) +
      (src04[60] << 4) +
      (src04[61] << 4) +
      (src04[62] << 4) +
      (src04[63] << 4) +
      (src05[0] << 5) +
      (src05[1] << 5) +
      (src05[2] << 5) +
      (src05[3] << 5) +
      (src05[4] << 5) +
      (src05[5] << 5) +
      (src05[6] << 5) +
      (src05[7] << 5) +
      (src05[8] << 5) +
      (src05[9] << 5) +
      (src05[10] << 5) +
      (src05[11] << 5) +
      (src05[12] << 5) +
      (src05[13] << 5) +
      (src05[14] << 5) +
      (src05[15] << 5) +
      (src05[16] << 5) +
      (src05[17] << 5) +
      (src05[18] << 5) +
      (src05[19] << 5) +
      (src05[20] << 5) +
      (src05[21] << 5) +
      (src05[22] << 5) +
      (src05[23] << 5) +
      (src05[24] << 5) +
      (src05[25] << 5) +
      (src05[26] << 5) +
      (src05[27] << 5) +
      (src05[28] << 5) +
      (src05[29] << 5) +
      (src05[30] << 5) +
      (src05[31] << 5) +
      (src05[32] << 5) +
      (src05[33] << 5) +
      (src05[34] << 5) +
      (src05[35] << 5) +
      (src05[36] << 5) +
      (src05[37] << 5) +
      (src05[38] << 5) +
      (src05[39] << 5) +
      (src05[40] << 5) +
      (src05[41] << 5) +
      (src05[42] << 5) +
      (src05[43] << 5) +
      (src05[44] << 5) +
      (src05[45] << 5) +
      (src05[46] << 5) +
      (src05[47] << 5) +
      (src05[48] << 5) +
      (src05[49] << 5) +
      (src05[50] << 5) +
      (src05[51] << 5) +
      (src05[52] << 5) +
      (src05[53] << 5) +
      (src05[54] << 5) +
      (src05[55] << 5) +
      (src05[56] << 5) +
      (src05[57] << 5) +
      (src05[58] << 5) +
      (src05[59] << 5) +
      (src05[60] << 5) +
      (src05[61] << 5) +
      (src05[62] << 5) +
      (src05[63] << 5) +
      (src06[0] << 6) +
      (src06[1] << 6) +
      (src06[2] << 6) +
      (src06[3] << 6) +
      (src06[4] << 6) +
      (src06[5] << 6) +
      (src06[6] << 6) +
      (src06[7] << 6) +
      (src06[8] << 6) +
      (src06[9] << 6) +
      (src06[10] << 6) +
      (src06[11] << 6) +
      (src06[12] << 6) +
      (src06[13] << 6) +
      (src06[14] << 6) +
      (src06[15] << 6) +
      (src06[16] << 6) +
      (src06[17] << 6) +
      (src06[18] << 6) +
      (src06[19] << 6) +
      (src06[20] << 6) +
      (src06[21] << 6) +
      (src06[22] << 6) +
      (src06[23] << 6) +
      (src06[24] << 6) +
      (src06[25] << 6) +
      (src06[26] << 6) +
      (src06[27] << 6) +
      (src06[28] << 6) +
      (src06[29] << 6) +
      (src06[30] << 6) +
      (src06[31] << 6) +
      (src06[32] << 6) +
      (src06[33] << 6) +
      (src06[34] << 6) +
      (src06[35] << 6) +
      (src06[36] << 6) +
      (src06[37] << 6) +
      (src06[38] << 6) +
      (src06[39] << 6) +
      (src06[40] << 6) +
      (src06[41] << 6) +
      (src06[42] << 6) +
      (src06[43] << 6) +
      (src06[44] << 6) +
      (src06[45] << 6) +
      (src06[46] << 6) +
      (src06[47] << 6) +
      (src06[48] << 6) +
      (src06[49] << 6) +
      (src06[50] << 6) +
      (src06[51] << 6) +
      (src06[52] << 6) +
      (src06[53] << 6) +
      (src06[54] << 6) +
      (src06[55] << 6) +
      (src06[56] << 6) +
      (src06[57] << 6) +
      (src06[58] << 6) +
      (src06[59] << 6) +
      (src06[60] << 6) +
      (src06[61] << 6) +
      (src06[62] << 6) +
      (src06[63] << 6) +
      (src07[0] << 7) +
      (src07[1] << 7) +
      (src07[2] << 7) +
      (src07[3] << 7) +
      (src07[4] << 7) +
      (src07[5] << 7) +
      (src07[6] << 7) +
      (src07[7] << 7) +
      (src07[8] << 7) +
      (src07[9] << 7) +
      (src07[10] << 7) +
      (src07[11] << 7) +
      (src07[12] << 7) +
      (src07[13] << 7) +
      (src07[14] << 7) +
      (src07[15] << 7) +
      (src07[16] << 7) +
      (src07[17] << 7) +
      (src07[18] << 7) +
      (src07[19] << 7) +
      (src07[20] << 7) +
      (src07[21] << 7) +
      (src07[22] << 7) +
      (src07[23] << 7) +
      (src07[24] << 7) +
      (src07[25] << 7) +
      (src07[26] << 7) +
      (src07[27] << 7) +
      (src07[28] << 7) +
      (src07[29] << 7) +
      (src07[30] << 7) +
      (src07[31] << 7) +
      (src07[32] << 7) +
      (src07[33] << 7) +
      (src07[34] << 7) +
      (src07[35] << 7) +
      (src07[36] << 7) +
      (src07[37] << 7) +
      (src07[38] << 7) +
      (src07[39] << 7) +
      (src07[40] << 7) +
      (src07[41] << 7) +
      (src07[42] << 7) +
      (src07[43] << 7) +
      (src07[44] << 7) +
      (src07[45] << 7) +
      (src07[46] << 7) +
      (src07[47] << 7) +
      (src07[48] << 7) +
      (src07[49] << 7) +
      (src07[50] << 7) +
      (src07[51] << 7) +
      (src07[52] << 7) +
      (src07[53] << 7) +
      (src07[54] << 7) +
      (src07[55] << 7) +
      (src07[56] << 7) +
      (src07[57] << 7) +
      (src07[58] << 7) +
      (src07[59] << 7) +
      (src07[60] << 7) +
      (src07[61] << 7) +
      (src07[62] << 7) +
      (src07[63] << 7) +
      (src08[0] << 8) +
      (src08[1] << 8) +
      (src08[2] << 8) +
      (src08[3] << 8) +
      (src08[4] << 8) +
      (src08[5] << 8) +
      (src08[6] << 8) +
      (src08[7] << 8) +
      (src08[8] << 8) +
      (src08[9] << 8) +
      (src08[10] << 8) +
      (src08[11] << 8) +
      (src08[12] << 8) +
      (src08[13] << 8) +
      (src08[14] << 8) +
      (src08[15] << 8) +
      (src08[16] << 8) +
      (src08[17] << 8) +
      (src08[18] << 8) +
      (src08[19] << 8) +
      (src08[20] << 8) +
      (src08[21] << 8) +
      (src08[22] << 8) +
      (src08[23] << 8) +
      (src08[24] << 8) +
      (src08[25] << 8) +
      (src08[26] << 8) +
      (src08[27] << 8) +
      (src08[28] << 8) +
      (src08[29] << 8) +
      (src08[30] << 8) +
      (src08[31] << 8) +
      (src08[32] << 8) +
      (src08[33] << 8) +
      (src08[34] << 8) +
      (src08[35] << 8) +
      (src08[36] << 8) +
      (src08[37] << 8) +
      (src08[38] << 8) +
      (src08[39] << 8) +
      (src08[40] << 8) +
      (src08[41] << 8) +
      (src08[42] << 8) +
      (src08[43] << 8) +
      (src08[44] << 8) +
      (src08[45] << 8) +
      (src08[46] << 8) +
      (src08[47] << 8) +
      (src08[48] << 8) +
      (src08[49] << 8) +
      (src08[50] << 8) +
      (src08[51] << 8) +
      (src08[52] << 8) +
      (src08[53] << 8) +
      (src08[54] << 8) +
      (src08[55] << 8) +
      (src08[56] << 8) +
      (src08[57] << 8) +
      (src08[58] << 8) +
      (src08[59] << 8) +
      (src08[60] << 8) +
      (src08[61] << 8) +
      (src08[62] << 8) +
      (src08[63] << 8) +
      (src09[0] << 9) +
      (src09[1] << 9) +
      (src09[2] << 9) +
      (src09[3] << 9) +
      (src09[4] << 9) +
      (src09[5] << 9) +
      (src09[6] << 9) +
      (src09[7] << 9) +
      (src09[8] << 9) +
      (src09[9] << 9) +
      (src09[10] << 9) +
      (src09[11] << 9) +
      (src09[12] << 9) +
      (src09[13] << 9) +
      (src09[14] << 9) +
      (src09[15] << 9) +
      (src09[16] << 9) +
      (src09[17] << 9) +
      (src09[18] << 9) +
      (src09[19] << 9) +
      (src09[20] << 9) +
      (src09[21] << 9) +
      (src09[22] << 9) +
      (src09[23] << 9) +
      (src09[24] << 9) +
      (src09[25] << 9) +
      (src09[26] << 9) +
      (src09[27] << 9) +
      (src09[28] << 9) +
      (src09[29] << 9) +
      (src09[30] << 9) +
      (src09[31] << 9) +
      (src09[32] << 9) +
      (src09[33] << 9) +
      (src09[34] << 9) +
      (src09[35] << 9) +
      (src09[36] << 9) +
      (src09[37] << 9) +
      (src09[38] << 9) +
      (src09[39] << 9) +
      (src09[40] << 9) +
      (src09[41] << 9) +
      (src09[42] << 9) +
      (src09[43] << 9) +
      (src09[44] << 9) +
      (src09[45] << 9) +
      (src09[46] << 9) +
      (src09[47] << 9) +
      (src09[48] << 9) +
      (src09[49] << 9) +
      (src09[50] << 9) +
      (src09[51] << 9) +
      (src09[52] << 9) +
      (src09[53] << 9) +
      (src09[54] << 9) +
      (src09[55] << 9) +
      (src09[56] << 9) +
      (src09[57] << 9) +
      (src09[58] << 9) +
      (src09[59] << 9) +
      (src09[60] << 9) +
      (src09[61] << 9) +
      (src09[62] << 9) +
      (src09[63] << 9) +
      (src10[0] << 10) +
      (src10[1] << 10) +
      (src10[2] << 10) +
      (src10[3] << 10) +
      (src10[4] << 10) +
      (src10[5] << 10) +
      (src10[6] << 10) +
      (src10[7] << 10) +
      (src10[8] << 10) +
      (src10[9] << 10) +
      (src10[10] << 10) +
      (src10[11] << 10) +
      (src10[12] << 10) +
      (src10[13] << 10) +
      (src10[14] << 10) +
      (src10[15] << 10) +
      (src10[16] << 10) +
      (src10[17] << 10) +
      (src10[18] << 10) +
      (src10[19] << 10) +
      (src10[20] << 10) +
      (src10[21] << 10) +
      (src10[22] << 10) +
      (src10[23] << 10) +
      (src10[24] << 10) +
      (src10[25] << 10) +
      (src10[26] << 10) +
      (src10[27] << 10) +
      (src10[28] << 10) +
      (src10[29] << 10) +
      (src10[30] << 10) +
      (src10[31] << 10) +
      (src10[32] << 10) +
      (src10[33] << 10) +
      (src10[34] << 10) +
      (src10[35] << 10) +
      (src10[36] << 10) +
      (src10[37] << 10) +
      (src10[38] << 10) +
      (src10[39] << 10) +
      (src10[40] << 10) +
      (src10[41] << 10) +
      (src10[42] << 10) +
      (src10[43] << 10) +
      (src10[44] << 10) +
      (src10[45] << 10) +
      (src10[46] << 10) +
      (src10[47] << 10) +
      (src10[48] << 10) +
      (src10[49] << 10) +
      (src10[50] << 10) +
      (src10[51] << 10) +
      (src10[52] << 10) +
      (src10[53] << 10) +
      (src10[54] << 10) +
      (src10[55] << 10) +
      (src10[56] << 10) +
      (src10[57] << 10) +
      (src10[58] << 10) +
      (src10[59] << 10) +
      (src10[60] << 10) +
      (src10[61] << 10) +
      (src10[62] << 10) +
      (src10[63] << 10) +
      (src11[0] << 11) +
      (src11[1] << 11) +
      (src11[2] << 11) +
      (src11[3] << 11) +
      (src11[4] << 11) +
      (src11[5] << 11) +
      (src11[6] << 11) +
      (src11[7] << 11) +
      (src11[8] << 11) +
      (src11[9] << 11) +
      (src11[10] << 11) +
      (src11[11] << 11) +
      (src11[12] << 11) +
      (src11[13] << 11) +
      (src11[14] << 11) +
      (src11[15] << 11) +
      (src11[16] << 11) +
      (src11[17] << 11) +
      (src11[18] << 11) +
      (src11[19] << 11) +
      (src11[20] << 11) +
      (src11[21] << 11) +
      (src11[22] << 11) +
      (src11[23] << 11) +
      (src11[24] << 11) +
      (src11[25] << 11) +
      (src11[26] << 11) +
      (src11[27] << 11) +
      (src11[28] << 11) +
      (src11[29] << 11) +
      (src11[30] << 11) +
      (src11[31] << 11) +
      (src11[32] << 11) +
      (src11[33] << 11) +
      (src11[34] << 11) +
      (src11[35] << 11) +
      (src11[36] << 11) +
      (src11[37] << 11) +
      (src11[38] << 11) +
      (src11[39] << 11) +
      (src11[40] << 11) +
      (src11[41] << 11) +
      (src11[42] << 11) +
      (src11[43] << 11) +
      (src11[44] << 11) +
      (src11[45] << 11) +
      (src11[46] << 11) +
      (src11[47] << 11) +
      (src11[48] << 11) +
      (src11[49] << 11) +
      (src11[50] << 11) +
      (src11[51] << 11) +
      (src11[52] << 11) +
      (src11[53] << 11) +
      (src11[54] << 11) +
      (src11[55] << 11) +
      (src11[56] << 11) +
      (src11[57] << 11) +
      (src11[58] << 11) +
      (src11[59] << 11) +
      (src11[60] << 11) +
      (src11[61] << 11) +
      (src11[62] << 11) +
      (src11[63] << 11) +
      (src12[0] << 12) +
      (src12[1] << 12) +
      (src12[2] << 12) +
      (src12[3] << 12) +
      (src12[4] << 12) +
      (src12[5] << 12) +
      (src12[6] << 12) +
      (src12[7] << 12) +
      (src12[8] << 12) +
      (src12[9] << 12) +
      (src12[10] << 12) +
      (src12[11] << 12) +
      (src12[12] << 12) +
      (src12[13] << 12) +
      (src12[14] << 12) +
      (src12[15] << 12) +
      (src12[16] << 12) +
      (src12[17] << 12) +
      (src12[18] << 12) +
      (src12[19] << 12) +
      (src12[20] << 12) +
      (src12[21] << 12) +
      (src12[22] << 12) +
      (src12[23] << 12) +
      (src12[24] << 12) +
      (src12[25] << 12) +
      (src12[26] << 12) +
      (src12[27] << 12) +
      (src12[28] << 12) +
      (src12[29] << 12) +
      (src12[30] << 12) +
      (src12[31] << 12) +
      (src12[32] << 12) +
      (src12[33] << 12) +
      (src12[34] << 12) +
      (src12[35] << 12) +
      (src12[36] << 12) +
      (src12[37] << 12) +
      (src12[38] << 12) +
      (src12[39] << 12) +
      (src12[40] << 12) +
      (src12[41] << 12) +
      (src12[42] << 12) +
      (src12[43] << 12) +
      (src12[44] << 12) +
      (src12[45] << 12) +
      (src12[46] << 12) +
      (src12[47] << 12) +
      (src12[48] << 12) +
      (src12[49] << 12) +
      (src12[50] << 12) +
      (src12[51] << 12) +
      (src12[52] << 12) +
      (src12[53] << 12) +
      (src12[54] << 12) +
      (src12[55] << 12) +
      (src12[56] << 12) +
      (src12[57] << 12) +
      (src12[58] << 12) +
      (src12[59] << 12) +
      (src12[60] << 12) +
      (src12[61] << 12) +
      (src12[62] << 12) +
      (src12[63] << 12) +
      (src13[0] << 13) +
      (src13[1] << 13) +
      (src13[2] << 13) +
      (src13[3] << 13) +
      (src13[4] << 13) +
      (src13[5] << 13) +
      (src13[6] << 13) +
      (src13[7] << 13) +
      (src13[8] << 13) +
      (src13[9] << 13) +
      (src13[10] << 13) +
      (src13[11] << 13) +
      (src13[12] << 13) +
      (src13[13] << 13) +
      (src13[14] << 13) +
      (src13[15] << 13) +
      (src13[16] << 13) +
      (src13[17] << 13) +
      (src13[18] << 13) +
      (src13[19] << 13) +
      (src13[20] << 13) +
      (src13[21] << 13) +
      (src13[22] << 13) +
      (src13[23] << 13) +
      (src13[24] << 13) +
      (src13[25] << 13) +
      (src13[26] << 13) +
      (src13[27] << 13) +
      (src13[28] << 13) +
      (src13[29] << 13) +
      (src13[30] << 13) +
      (src13[31] << 13) +
      (src13[32] << 13) +
      (src13[33] << 13) +
      (src13[34] << 13) +
      (src13[35] << 13) +
      (src13[36] << 13) +
      (src13[37] << 13) +
      (src13[38] << 13) +
      (src13[39] << 13) +
      (src13[40] << 13) +
      (src13[41] << 13) +
      (src13[42] << 13) +
      (src13[43] << 13) +
      (src13[44] << 13) +
      (src13[45] << 13) +
      (src13[46] << 13) +
      (src13[47] << 13) +
      (src13[48] << 13) +
      (src13[49] << 13) +
      (src13[50] << 13) +
      (src13[51] << 13) +
      (src13[52] << 13) +
      (src13[53] << 13) +
      (src13[54] << 13) +
      (src13[55] << 13) +
      (src13[56] << 13) +
      (src13[57] << 13) +
      (src13[58] << 13) +
      (src13[59] << 13) +
      (src13[60] << 13) +
      (src13[61] << 13) +
      (src13[62] << 13) +
      (src13[63] << 13) +
      (src14[0] << 14) +
      (src14[1] << 14) +
      (src14[2] << 14) +
      (src14[3] << 14) +
      (src14[4] << 14) +
      (src14[5] << 14) +
      (src14[6] << 14) +
      (src14[7] << 14) +
      (src14[8] << 14) +
      (src14[9] << 14) +
      (src14[10] << 14) +
      (src14[11] << 14) +
      (src14[12] << 14) +
      (src14[13] << 14) +
      (src14[14] << 14) +
      (src14[15] << 14) +
      (src14[16] << 14) +
      (src14[17] << 14) +
      (src14[18] << 14) +
      (src14[19] << 14) +
      (src14[20] << 14) +
      (src14[21] << 14) +
      (src14[22] << 14) +
      (src14[23] << 14) +
      (src14[24] << 14) +
      (src14[25] << 14) +
      (src14[26] << 14) +
      (src14[27] << 14) +
      (src14[28] << 14) +
      (src14[29] << 14) +
      (src14[30] << 14) +
      (src14[31] << 14) +
      (src14[32] << 14) +
      (src14[33] << 14) +
      (src14[34] << 14) +
      (src14[35] << 14) +
      (src14[36] << 14) +
      (src14[37] << 14) +
      (src14[38] << 14) +
      (src14[39] << 14) +
      (src14[40] << 14) +
      (src14[41] << 14) +
      (src14[42] << 14) +
      (src14[43] << 14) +
      (src14[44] << 14) +
      (src14[45] << 14) +
      (src14[46] << 14) +
      (src14[47] << 14) +
      (src14[48] << 14) +
      (src14[49] << 14) +
      (src14[50] << 14) +
      (src14[51] << 14) +
      (src14[52] << 14) +
      (src14[53] << 14) +
      (src14[54] << 14) +
      (src14[55] << 14) +
      (src14[56] << 14) +
      (src14[57] << 14) +
      (src14[58] << 14) +
      (src14[59] << 14) +
      (src14[60] << 14) +
      (src14[61] << 14) +
      (src14[62] << 14) +
      (src14[63] << 14) +
      (src15[0] << 15) +
      (src15[1] << 15) +
      (src15[2] << 15) +
      (src15[3] << 15) +
      (src15[4] << 15) +
      (src15[5] << 15) +
      (src15[6] << 15) +
      (src15[7] << 15) +
      (src15[8] << 15) +
      (src15[9] << 15) +
      (src15[10] << 15) +
      (src15[11] << 15) +
      (src15[12] << 15) +
      (src15[13] << 15) +
      (src15[14] << 15) +
      (src15[15] << 15) +
      (src15[16] << 15) +
      (src15[17] << 15) +
      (src15[18] << 15) +
      (src15[19] << 15) +
      (src15[20] << 15) +
      (src15[21] << 15) +
      (src15[22] << 15) +
      (src15[23] << 15) +
      (src15[24] << 15) +
      (src15[25] << 15) +
      (src15[26] << 15) +
      (src15[27] << 15) +
      (src15[28] << 15) +
      (src15[29] << 15) +
      (src15[30] << 15) +
      (src15[31] << 15) +
      (src15[32] << 15) +
      (src15[33] << 15) +
      (src15[34] << 15) +
      (src15[35] << 15) +
      (src15[36] << 15) +
      (src15[37] << 15) +
      (src15[38] << 15) +
      (src15[39] << 15) +
      (src15[40] << 15) +
      (src15[41] << 15) +
      (src15[42] << 15) +
      (src15[43] << 15) +
      (src15[44] << 15) +
      (src15[45] << 15) +
      (src15[46] << 15) +
      (src15[47] << 15) +
      (src15[48] << 15) +
      (src15[49] << 15) +
      (src15[50] << 15) +
      (src15[51] << 15) +
      (src15[52] << 15) +
      (src15[53] << 15) +
      (src15[54] << 15) +
      (src15[55] << 15) +
      (src15[56] << 15) +
      (src15[57] << 15) +
      (src15[58] << 15) +
      (src15[59] << 15) +
      (src15[60] << 15) +
      (src15[61] << 15) +
      (src15[62] << 15) +
      (src15[63] << 15) +
      (src16[0] << 16) +
      (src16[1] << 16) +
      (src16[2] << 16) +
      (src16[3] << 16) +
      (src16[4] << 16) +
      (src16[5] << 16) +
      (src16[6] << 16) +
      (src16[7] << 16) +
      (src16[8] << 16) +
      (src16[9] << 16) +
      (src16[10] << 16) +
      (src16[11] << 16) +
      (src16[12] << 16) +
      (src16[13] << 16) +
      (src16[14] << 16) +
      (src16[15] << 16) +
      (src16[16] << 16) +
      (src16[17] << 16) +
      (src16[18] << 16) +
      (src16[19] << 16) +
      (src16[20] << 16) +
      (src16[21] << 16) +
      (src16[22] << 16) +
      (src16[23] << 16) +
      (src16[24] << 16) +
      (src16[25] << 16) +
      (src16[26] << 16) +
      (src16[27] << 16) +
      (src16[28] << 16) +
      (src16[29] << 16) +
      (src16[30] << 16) +
      (src16[31] << 16) +
      (src16[32] << 16) +
      (src16[33] << 16) +
      (src16[34] << 16) +
      (src16[35] << 16) +
      (src16[36] << 16) +
      (src16[37] << 16) +
      (src16[38] << 16) +
      (src16[39] << 16) +
      (src16[40] << 16) +
      (src16[41] << 16) +
      (src16[42] << 16) +
      (src16[43] << 16) +
      (src16[44] << 16) +
      (src16[45] << 16) +
      (src16[46] << 16) +
      (src16[47] << 16) +
      (src16[48] << 16) +
      (src16[49] << 16) +
      (src16[50] << 16) +
      (src16[51] << 16) +
      (src16[52] << 16) +
      (src16[53] << 16) +
      (src16[54] << 16) +
      (src16[55] << 16) +
      (src16[56] << 16) +
      (src16[57] << 16) +
      (src16[58] << 16) +
      (src16[59] << 16) +
      (src16[60] << 16) +
      (src16[61] << 16) +
      (src16[62] << 16) +
      (src16[63] << 16) +
      (src17[0] << 17) +
      (src17[1] << 17) +
      (src17[2] << 17) +
      (src17[3] << 17) +
      (src17[4] << 17) +
      (src17[5] << 17) +
      (src17[6] << 17) +
      (src17[7] << 17) +
      (src17[8] << 17) +
      (src17[9] << 17) +
      (src17[10] << 17) +
      (src17[11] << 17) +
      (src17[12] << 17) +
      (src17[13] << 17) +
      (src17[14] << 17) +
      (src17[15] << 17) +
      (src17[16] << 17) +
      (src17[17] << 17) +
      (src17[18] << 17) +
      (src17[19] << 17) +
      (src17[20] << 17) +
      (src17[21] << 17) +
      (src17[22] << 17) +
      (src17[23] << 17) +
      (src17[24] << 17) +
      (src17[25] << 17) +
      (src17[26] << 17) +
      (src17[27] << 17) +
      (src17[28] << 17) +
      (src17[29] << 17) +
      (src17[30] << 17) +
      (src17[31] << 17) +
      (src17[32] << 17) +
      (src17[33] << 17) +
      (src17[34] << 17) +
      (src17[35] << 17) +
      (src17[36] << 17) +
      (src17[37] << 17) +
      (src17[38] << 17) +
      (src17[39] << 17) +
      (src17[40] << 17) +
      (src17[41] << 17) +
      (src17[42] << 17) +
      (src17[43] << 17) +
      (src17[44] << 17) +
      (src17[45] << 17) +
      (src17[46] << 17) +
      (src17[47] << 17) +
      (src17[48] << 17) +
      (src17[49] << 17) +
      (src17[50] << 17) +
      (src17[51] << 17) +
      (src17[52] << 17) +
      (src17[53] << 17) +
      (src17[54] << 17) +
      (src17[55] << 17) +
      (src17[56] << 17) +
      (src17[57] << 17) +
      (src17[58] << 17) +
      (src17[59] << 17) +
      (src17[60] << 17) +
      (src17[61] << 17) +
      (src17[62] << 17) +
      (src17[63] << 17) +
      (src18[0] << 18) +
      (src18[1] << 18) +
      (src18[2] << 18) +
      (src18[3] << 18) +
      (src18[4] << 18) +
      (src18[5] << 18) +
      (src18[6] << 18) +
      (src18[7] << 18) +
      (src18[8] << 18) +
      (src18[9] << 18) +
      (src18[10] << 18) +
      (src18[11] << 18) +
      (src18[12] << 18) +
      (src18[13] << 18) +
      (src18[14] << 18) +
      (src18[15] << 18) +
      (src18[16] << 18) +
      (src18[17] << 18) +
      (src18[18] << 18) +
      (src18[19] << 18) +
      (src18[20] << 18) +
      (src18[21] << 18) +
      (src18[22] << 18) +
      (src18[23] << 18) +
      (src18[24] << 18) +
      (src18[25] << 18) +
      (src18[26] << 18) +
      (src18[27] << 18) +
      (src18[28] << 18) +
      (src18[29] << 18) +
      (src18[30] << 18) +
      (src18[31] << 18) +
      (src18[32] << 18) +
      (src18[33] << 18) +
      (src18[34] << 18) +
      (src18[35] << 18) +
      (src18[36] << 18) +
      (src18[37] << 18) +
      (src18[38] << 18) +
      (src18[39] << 18) +
      (src18[40] << 18) +
      (src18[41] << 18) +
      (src18[42] << 18) +
      (src18[43] << 18) +
      (src18[44] << 18) +
      (src18[45] << 18) +
      (src18[46] << 18) +
      (src18[47] << 18) +
      (src18[48] << 18) +
      (src18[49] << 18) +
      (src18[50] << 18) +
      (src18[51] << 18) +
      (src18[52] << 18) +
      (src18[53] << 18) +
      (src18[54] << 18) +
      (src18[55] << 18) +
      (src18[56] << 18) +
      (src18[57] << 18) +
      (src18[58] << 18) +
      (src18[59] << 18) +
      (src18[60] << 18) +
      (src18[61] << 18) +
      (src18[62] << 18) +
      (src18[63] << 18) +
      (src19[0] << 19) +
      (src19[1] << 19) +
      (src19[2] << 19) +
      (src19[3] << 19) +
      (src19[4] << 19) +
      (src19[5] << 19) +
      (src19[6] << 19) +
      (src19[7] << 19) +
      (src19[8] << 19) +
      (src19[9] << 19) +
      (src19[10] << 19) +
      (src19[11] << 19) +
      (src19[12] << 19) +
      (src19[13] << 19) +
      (src19[14] << 19) +
      (src19[15] << 19) +
      (src19[16] << 19) +
      (src19[17] << 19) +
      (src19[18] << 19) +
      (src19[19] << 19) +
      (src19[20] << 19) +
      (src19[21] << 19) +
      (src19[22] << 19) +
      (src19[23] << 19) +
      (src19[24] << 19) +
      (src19[25] << 19) +
      (src19[26] << 19) +
      (src19[27] << 19) +
      (src19[28] << 19) +
      (src19[29] << 19) +
      (src19[30] << 19) +
      (src19[31] << 19) +
      (src19[32] << 19) +
      (src19[33] << 19) +
      (src19[34] << 19) +
      (src19[35] << 19) +
      (src19[36] << 19) +
      (src19[37] << 19) +
      (src19[38] << 19) +
      (src19[39] << 19) +
      (src19[40] << 19) +
      (src19[41] << 19) +
      (src19[42] << 19) +
      (src19[43] << 19) +
      (src19[44] << 19) +
      (src19[45] << 19) +
      (src19[46] << 19) +
      (src19[47] << 19) +
      (src19[48] << 19) +
      (src19[49] << 19) +
      (src19[50] << 19) +
      (src19[51] << 19) +
      (src19[52] << 19) +
      (src19[53] << 19) +
      (src19[54] << 19) +
      (src19[55] << 19) +
      (src19[56] << 19) +
      (src19[57] << 19) +
      (src19[58] << 19) +
      (src19[59] << 19) +
      (src19[60] << 19) +
      (src19[61] << 19) +
      (src19[62] << 19) +
      (src19[63] << 19) +
      (src20[0] << 20) +
      (src20[1] << 20) +
      (src20[2] << 20) +
      (src20[3] << 20) +
      (src20[4] << 20) +
      (src20[5] << 20) +
      (src20[6] << 20) +
      (src20[7] << 20) +
      (src20[8] << 20) +
      (src20[9] << 20) +
      (src20[10] << 20) +
      (src20[11] << 20) +
      (src20[12] << 20) +
      (src20[13] << 20) +
      (src20[14] << 20) +
      (src20[15] << 20) +
      (src20[16] << 20) +
      (src20[17] << 20) +
      (src20[18] << 20) +
      (src20[19] << 20) +
      (src20[20] << 20) +
      (src20[21] << 20) +
      (src20[22] << 20) +
      (src20[23] << 20) +
      (src20[24] << 20) +
      (src20[25] << 20) +
      (src20[26] << 20) +
      (src20[27] << 20) +
      (src20[28] << 20) +
      (src20[29] << 20) +
      (src20[30] << 20) +
      (src20[31] << 20) +
      (src20[32] << 20) +
      (src20[33] << 20) +
      (src20[34] << 20) +
      (src20[35] << 20) +
      (src20[36] << 20) +
      (src20[37] << 20) +
      (src20[38] << 20) +
      (src20[39] << 20) +
      (src20[40] << 20) +
      (src20[41] << 20) +
      (src20[42] << 20) +
      (src20[43] << 20) +
      (src20[44] << 20) +
      (src20[45] << 20) +
      (src20[46] << 20) +
      (src20[47] << 20) +
      (src20[48] << 20) +
      (src20[49] << 20) +
      (src20[50] << 20) +
      (src20[51] << 20) +
      (src20[52] << 20) +
      (src20[53] << 20) +
      (src20[54] << 20) +
      (src20[55] << 20) +
      (src20[56] << 20) +
      (src20[57] << 20) +
      (src20[58] << 20) +
      (src20[59] << 20) +
      (src20[60] << 20) +
      (src20[61] << 20) +
      (src20[62] << 20) +
      (src20[63] << 20) +
      (src21[0] << 21) +
      (src21[1] << 21) +
      (src21[2] << 21) +
      (src21[3] << 21) +
      (src21[4] << 21) +
      (src21[5] << 21) +
      (src21[6] << 21) +
      (src21[7] << 21) +
      (src21[8] << 21) +
      (src21[9] << 21) +
      (src21[10] << 21) +
      (src21[11] << 21) +
      (src21[12] << 21) +
      (src21[13] << 21) +
      (src21[14] << 21) +
      (src21[15] << 21) +
      (src21[16] << 21) +
      (src21[17] << 21) +
      (src21[18] << 21) +
      (src21[19] << 21) +
      (src21[20] << 21) +
      (src21[21] << 21) +
      (src21[22] << 21) +
      (src21[23] << 21) +
      (src21[24] << 21) +
      (src21[25] << 21) +
      (src21[26] << 21) +
      (src21[27] << 21) +
      (src21[28] << 21) +
      (src21[29] << 21) +
      (src21[30] << 21) +
      (src21[31] << 21) +
      (src21[32] << 21) +
      (src21[33] << 21) +
      (src21[34] << 21) +
      (src21[35] << 21) +
      (src21[36] << 21) +
      (src21[37] << 21) +
      (src21[38] << 21) +
      (src21[39] << 21) +
      (src21[40] << 21) +
      (src21[41] << 21) +
      (src21[42] << 21) +
      (src21[43] << 21) +
      (src21[44] << 21) +
      (src21[45] << 21) +
      (src21[46] << 21) +
      (src21[47] << 21) +
      (src21[48] << 21) +
      (src21[49] << 21) +
      (src21[50] << 21) +
      (src21[51] << 21) +
      (src21[52] << 21) +
      (src21[53] << 21) +
      (src21[54] << 21) +
      (src21[55] << 21) +
      (src21[56] << 21) +
      (src21[57] << 21) +
      (src21[58] << 21) +
      (src21[59] << 21) +
      (src21[60] << 21) +
      (src21[61] << 21) +
      (src21[62] << 21) +
      (src21[63] << 21) +
      (src22[0] << 22) +
      (src22[1] << 22) +
      (src22[2] << 22) +
      (src22[3] << 22) +
      (src22[4] << 22) +
      (src22[5] << 22) +
      (src22[6] << 22) +
      (src22[7] << 22) +
      (src22[8] << 22) +
      (src22[9] << 22) +
      (src22[10] << 22) +
      (src22[11] << 22) +
      (src22[12] << 22) +
      (src22[13] << 22) +
      (src22[14] << 22) +
      (src22[15] << 22) +
      (src22[16] << 22) +
      (src22[17] << 22) +
      (src22[18] << 22) +
      (src22[19] << 22) +
      (src22[20] << 22) +
      (src22[21] << 22) +
      (src22[22] << 22) +
      (src22[23] << 22) +
      (src22[24] << 22) +
      (src22[25] << 22) +
      (src22[26] << 22) +
      (src22[27] << 22) +
      (src22[28] << 22) +
      (src22[29] << 22) +
      (src22[30] << 22) +
      (src22[31] << 22) +
      (src22[32] << 22) +
      (src22[33] << 22) +
      (src22[34] << 22) +
      (src22[35] << 22) +
      (src22[36] << 22) +
      (src22[37] << 22) +
      (src22[38] << 22) +
      (src22[39] << 22) +
      (src22[40] << 22) +
      (src22[41] << 22) +
      (src22[42] << 22) +
      (src22[43] << 22) +
      (src22[44] << 22) +
      (src22[45] << 22) +
      (src22[46] << 22) +
      (src22[47] << 22) +
      (src22[48] << 22) +
      (src22[49] << 22) +
      (src22[50] << 22) +
      (src22[51] << 22) +
      (src22[52] << 22) +
      (src22[53] << 22) +
      (src22[54] << 22) +
      (src22[55] << 22) +
      (src22[56] << 22) +
      (src22[57] << 22) +
      (src22[58] << 22) +
      (src22[59] << 22) +
      (src22[60] << 22) +
      (src22[61] << 22) +
      (src22[62] << 22) +
      (src22[63] << 22) +
      (src23[0] << 23) +
      (src23[1] << 23) +
      (src23[2] << 23) +
      (src23[3] << 23) +
      (src23[4] << 23) +
      (src23[5] << 23) +
      (src23[6] << 23) +
      (src23[7] << 23) +
      (src23[8] << 23) +
      (src23[9] << 23) +
      (src23[10] << 23) +
      (src23[11] << 23) +
      (src23[12] << 23) +
      (src23[13] << 23) +
      (src23[14] << 23) +
      (src23[15] << 23) +
      (src23[16] << 23) +
      (src23[17] << 23) +
      (src23[18] << 23) +
      (src23[19] << 23) +
      (src23[20] << 23) +
      (src23[21] << 23) +
      (src23[22] << 23) +
      (src23[23] << 23) +
      (src23[24] << 23) +
      (src23[25] << 23) +
      (src23[26] << 23) +
      (src23[27] << 23) +
      (src23[28] << 23) +
      (src23[29] << 23) +
      (src23[30] << 23) +
      (src23[31] << 23) +
      (src23[32] << 23) +
      (src23[33] << 23) +
      (src23[34] << 23) +
      (src23[35] << 23) +
      (src23[36] << 23) +
      (src23[37] << 23) +
      (src23[38] << 23) +
      (src23[39] << 23) +
      (src23[40] << 23) +
      (src23[41] << 23) +
      (src23[42] << 23) +
      (src23[43] << 23) +
      (src23[44] << 23) +
      (src23[45] << 23) +
      (src23[46] << 23) +
      (src23[47] << 23) +
      (src23[48] << 23) +
      (src23[49] << 23) +
      (src23[50] << 23) +
      (src23[51] << 23) +
      (src23[52] << 23) +
      (src23[53] << 23) +
      (src23[54] << 23) +
      (src23[55] << 23) +
      (src23[56] << 23) +
      (src23[57] << 23) +
      (src23[58] << 23) +
      (src23[59] << 23) +
      (src23[60] << 23) +
      (src23[61] << 23) +
      (src23[62] << 23) +
      (src23[63] << 23) +
      (src24[0] << 24) +
      (src24[1] << 24) +
      (src24[2] << 24) +
      (src24[3] << 24) +
      (src24[4] << 24) +
      (src24[5] << 24) +
      (src24[6] << 24) +
      (src24[7] << 24) +
      (src24[8] << 24) +
      (src24[9] << 24) +
      (src24[10] << 24) +
      (src24[11] << 24) +
      (src24[12] << 24) +
      (src24[13] << 24) +
      (src24[14] << 24) +
      (src24[15] << 24) +
      (src24[16] << 24) +
      (src24[17] << 24) +
      (src24[18] << 24) +
      (src24[19] << 24) +
      (src24[20] << 24) +
      (src24[21] << 24) +
      (src24[22] << 24) +
      (src24[23] << 24) +
      (src24[24] << 24) +
      (src24[25] << 24) +
      (src24[26] << 24) +
      (src24[27] << 24) +
      (src24[28] << 24) +
      (src24[29] << 24) +
      (src24[30] << 24) +
      (src24[31] << 24) +
      (src24[32] << 24) +
      (src24[33] << 24) +
      (src24[34] << 24) +
      (src24[35] << 24) +
      (src24[36] << 24) +
      (src24[37] << 24) +
      (src24[38] << 24) +
      (src24[39] << 24) +
      (src24[40] << 24) +
      (src24[41] << 24) +
      (src24[42] << 24) +
      (src24[43] << 24) +
      (src24[44] << 24) +
      (src24[45] << 24) +
      (src24[46] << 24) +
      (src24[47] << 24) +
      (src24[48] << 24) +
      (src24[49] << 24) +
      (src24[50] << 24) +
      (src24[51] << 24) +
      (src24[52] << 24) +
      (src24[53] << 24) +
      (src24[54] << 24) +
      (src24[55] << 24) +
      (src24[56] << 24) +
      (src24[57] << 24) +
      (src24[58] << 24) +
      (src24[59] << 24) +
      (src24[60] << 24) +
      (src24[61] << 24) +
      (src24[62] << 24) +
      (src24[63] << 24) +
      (src25[0] << 25) +
      (src25[1] << 25) +
      (src25[2] << 25) +
      (src25[3] << 25) +
      (src25[4] << 25) +
      (src25[5] << 25) +
      (src25[6] << 25) +
      (src25[7] << 25) +
      (src25[8] << 25) +
      (src25[9] << 25) +
      (src25[10] << 25) +
      (src25[11] << 25) +
      (src25[12] << 25) +
      (src25[13] << 25) +
      (src25[14] << 25) +
      (src25[15] << 25) +
      (src25[16] << 25) +
      (src25[17] << 25) +
      (src25[18] << 25) +
      (src25[19] << 25) +
      (src25[20] << 25) +
      (src25[21] << 25) +
      (src25[22] << 25) +
      (src25[23] << 25) +
      (src25[24] << 25) +
      (src25[25] << 25) +
      (src25[26] << 25) +
      (src25[27] << 25) +
      (src25[28] << 25) +
      (src25[29] << 25) +
      (src25[30] << 25) +
      (src25[31] << 25) +
      (src25[32] << 25) +
      (src25[33] << 25) +
      (src25[34] << 25) +
      (src25[35] << 25) +
      (src25[36] << 25) +
      (src25[37] << 25) +
      (src25[38] << 25) +
      (src25[39] << 25) +
      (src25[40] << 25) +
      (src25[41] << 25) +
      (src25[42] << 25) +
      (src25[43] << 25) +
      (src25[44] << 25) +
      (src25[45] << 25) +
      (src25[46] << 25) +
      (src25[47] << 25) +
      (src25[48] << 25) +
      (src25[49] << 25) +
      (src25[50] << 25) +
      (src25[51] << 25) +
      (src25[52] << 25) +
      (src25[53] << 25) +
      (src25[54] << 25) +
      (src25[55] << 25) +
      (src25[56] << 25) +
      (src25[57] << 25) +
      (src25[58] << 25) +
      (src25[59] << 25) +
      (src25[60] << 25) +
      (src25[61] << 25) +
      (src25[62] << 25) +
      (src25[63] << 25) +
      (src26[0] << 26) +
      (src26[1] << 26) +
      (src26[2] << 26) +
      (src26[3] << 26) +
      (src26[4] << 26) +
      (src26[5] << 26) +
      (src26[6] << 26) +
      (src26[7] << 26) +
      (src26[8] << 26) +
      (src26[9] << 26) +
      (src26[10] << 26) +
      (src26[11] << 26) +
      (src26[12] << 26) +
      (src26[13] << 26) +
      (src26[14] << 26) +
      (src26[15] << 26) +
      (src26[16] << 26) +
      (src26[17] << 26) +
      (src26[18] << 26) +
      (src26[19] << 26) +
      (src26[20] << 26) +
      (src26[21] << 26) +
      (src26[22] << 26) +
      (src26[23] << 26) +
      (src26[24] << 26) +
      (src26[25] << 26) +
      (src26[26] << 26) +
      (src26[27] << 26) +
      (src26[28] << 26) +
      (src26[29] << 26) +
      (src26[30] << 26) +
      (src26[31] << 26) +
      (src26[32] << 26) +
      (src26[33] << 26) +
      (src26[34] << 26) +
      (src26[35] << 26) +
      (src26[36] << 26) +
      (src26[37] << 26) +
      (src26[38] << 26) +
      (src26[39] << 26) +
      (src26[40] << 26) +
      (src26[41] << 26) +
      (src26[42] << 26) +
      (src26[43] << 26) +
      (src26[44] << 26) +
      (src26[45] << 26) +
      (src26[46] << 26) +
      (src26[47] << 26) +
      (src26[48] << 26) +
      (src26[49] << 26) +
      (src26[50] << 26) +
      (src26[51] << 26) +
      (src26[52] << 26) +
      (src26[53] << 26) +
      (src26[54] << 26) +
      (src26[55] << 26) +
      (src26[56] << 26) +
      (src26[57] << 26) +
      (src26[58] << 26) +
      (src26[59] << 26) +
      (src26[60] << 26) +
      (src26[61] << 26) +
      (src26[62] << 26) +
      (src26[63] << 26) +
      (src27[0] << 27) +
      (src27[1] << 27) +
      (src27[2] << 27) +
      (src27[3] << 27) +
      (src27[4] << 27) +
      (src27[5] << 27) +
      (src27[6] << 27) +
      (src27[7] << 27) +
      (src27[8] << 27) +
      (src27[9] << 27) +
      (src27[10] << 27) +
      (src27[11] << 27) +
      (src27[12] << 27) +
      (src27[13] << 27) +
      (src27[14] << 27) +
      (src27[15] << 27) +
      (src27[16] << 27) +
      (src27[17] << 27) +
      (src27[18] << 27) +
      (src27[19] << 27) +
      (src27[20] << 27) +
      (src27[21] << 27) +
      (src27[22] << 27) +
      (src27[23] << 27) +
      (src27[24] << 27) +
      (src27[25] << 27) +
      (src27[26] << 27) +
      (src27[27] << 27) +
      (src27[28] << 27) +
      (src27[29] << 27) +
      (src27[30] << 27) +
      (src27[31] << 27) +
      (src27[32] << 27) +
      (src27[33] << 27) +
      (src27[34] << 27) +
      (src27[35] << 27) +
      (src27[36] << 27) +
      (src27[37] << 27) +
      (src27[38] << 27) +
      (src27[39] << 27) +
      (src27[40] << 27) +
      (src27[41] << 27) +
      (src27[42] << 27) +
      (src27[43] << 27) +
      (src27[44] << 27) +
      (src27[45] << 27) +
      (src27[46] << 27) +
      (src27[47] << 27) +
      (src27[48] << 27) +
      (src27[49] << 27) +
      (src27[50] << 27) +
      (src27[51] << 27) +
      (src27[52] << 27) +
      (src27[53] << 27) +
      (src27[54] << 27) +
      (src27[55] << 27) +
      (src27[56] << 27) +
      (src27[57] << 27) +
      (src27[58] << 27) +
      (src27[59] << 27) +
      (src27[60] << 27) +
      (src27[61] << 27) +
      (src27[62] << 27) +
      (src27[63] << 27) +
      (src28[0] << 28) +
      (src28[1] << 28) +
      (src28[2] << 28) +
      (src28[3] << 28) +
      (src28[4] << 28) +
      (src28[5] << 28) +
      (src28[6] << 28) +
      (src28[7] << 28) +
      (src28[8] << 28) +
      (src28[9] << 28) +
      (src28[10] << 28) +
      (src28[11] << 28) +
      (src28[12] << 28) +
      (src28[13] << 28) +
      (src28[14] << 28) +
      (src28[15] << 28) +
      (src28[16] << 28) +
      (src28[17] << 28) +
      (src28[18] << 28) +
      (src28[19] << 28) +
      (src28[20] << 28) +
      (src28[21] << 28) +
      (src28[22] << 28) +
      (src28[23] << 28) +
      (src28[24] << 28) +
      (src28[25] << 28) +
      (src28[26] << 28) +
      (src28[27] << 28) +
      (src28[28] << 28) +
      (src28[29] << 28) +
      (src28[30] << 28) +
      (src28[31] << 28) +
      (src28[32] << 28) +
      (src28[33] << 28) +
      (src28[34] << 28) +
      (src28[35] << 28) +
      (src28[36] << 28) +
      (src28[37] << 28) +
      (src28[38] << 28) +
      (src28[39] << 28) +
      (src28[40] << 28) +
      (src28[41] << 28) +
      (src28[42] << 28) +
      (src28[43] << 28) +
      (src28[44] << 28) +
      (src28[45] << 28) +
      (src28[46] << 28) +
      (src28[47] << 28) +
      (src28[48] << 28) +
      (src28[49] << 28) +
      (src28[50] << 28) +
      (src28[51] << 28) +
      (src28[52] << 28) +
      (src28[53] << 28) +
      (src28[54] << 28) +
      (src28[55] << 28) +
      (src28[56] << 28) +
      (src28[57] << 28) +
      (src28[58] << 28) +
      (src28[59] << 28) +
      (src28[60] << 28) +
      (src28[61] << 28) +
      (src28[62] << 28) +
      (src28[63] << 28) +
      (src29[0] << 29) +
      (src29[1] << 29) +
      (src29[2] << 29) +
      (src29[3] << 29) +
      (src29[4] << 29) +
      (src29[5] << 29) +
      (src29[6] << 29) +
      (src29[7] << 29) +
      (src29[8] << 29) +
      (src29[9] << 29) +
      (src29[10] << 29) +
      (src29[11] << 29) +
      (src29[12] << 29) +
      (src29[13] << 29) +
      (src29[14] << 29) +
      (src29[15] << 29) +
      (src29[16] << 29) +
      (src29[17] << 29) +
      (src29[18] << 29) +
      (src29[19] << 29) +
      (src29[20] << 29) +
      (src29[21] << 29) +
      (src29[22] << 29) +
      (src29[23] << 29) +
      (src29[24] << 29) +
      (src29[25] << 29) +
      (src29[26] << 29) +
      (src29[27] << 29) +
      (src29[28] << 29) +
      (src29[29] << 29) +
      (src29[30] << 29) +
      (src29[31] << 29) +
      (src29[32] << 29) +
      (src29[33] << 29) +
      (src29[34] << 29) +
      (src29[35] << 29) +
      (src29[36] << 29) +
      (src29[37] << 29) +
      (src29[38] << 29) +
      (src29[39] << 29) +
      (src29[40] << 29) +
      (src29[41] << 29) +
      (src29[42] << 29) +
      (src29[43] << 29) +
      (src29[44] << 29) +
      (src29[45] << 29) +
      (src29[46] << 29) +
      (src29[47] << 29) +
      (src29[48] << 29) +
      (src29[49] << 29) +
      (src29[50] << 29) +
      (src29[51] << 29) +
      (src29[52] << 29) +
      (src29[53] << 29) +
      (src29[54] << 29) +
      (src29[55] << 29) +
      (src29[56] << 29) +
      (src29[57] << 29) +
      (src29[58] << 29) +
      (src29[59] << 29) +
      (src29[60] << 29) +
      (src29[61] << 29) +
      (src29[62] << 29) +
      (src29[63] << 29) +
      (src30[0] << 30) +
      (src30[1] << 30) +
      (src30[2] << 30) +
      (src30[3] << 30) +
      (src30[4] << 30) +
      (src30[5] << 30) +
      (src30[6] << 30) +
      (src30[7] << 30) +
      (src30[8] << 30) +
      (src30[9] << 30) +
      (src30[10] << 30) +
      (src30[11] << 30) +
      (src30[12] << 30) +
      (src30[13] << 30) +
      (src30[14] << 30) +
      (src30[15] << 30) +
      (src30[16] << 30) +
      (src30[17] << 30) +
      (src30[18] << 30) +
      (src30[19] << 30) +
      (src30[20] << 30) +
      (src30[21] << 30) +
      (src30[22] << 30) +
      (src30[23] << 30) +
      (src30[24] << 30) +
      (src30[25] << 30) +
      (src30[26] << 30) +
      (src30[27] << 30) +
      (src30[28] << 30) +
      (src30[29] << 30) +
      (src30[30] << 30) +
      (src30[31] << 30) +
      (src30[32] << 30) +
      (src30[33] << 30) +
      (src30[34] << 30) +
      (src30[35] << 30) +
      (src30[36] << 30) +
      (src30[37] << 30) +
      (src30[38] << 30) +
      (src30[39] << 30) +
      (src30[40] << 30) +
      (src30[41] << 30) +
      (src30[42] << 30) +
      (src30[43] << 30) +
      (src30[44] << 30) +
      (src30[45] << 30) +
      (src30[46] << 30) +
      (src30[47] << 30) +
      (src30[48] << 30) +
      (src30[49] << 30) +
      (src30[50] << 30) +
      (src30[51] << 30) +
      (src30[52] << 30) +
      (src30[53] << 30) +
      (src30[54] << 30) +
      (src30[55] << 30) +
      (src30[56] << 30) +
      (src30[57] << 30) +
      (src30[58] << 30) +
      (src30[59] << 30) +
      (src30[60] << 30) +
      (src30[61] << 30) +
      (src30[62] << 30) +
      (src30[63] << 30) +
      (src31[0] << 31) +
      (src31[1] << 31) +
      (src31[2] << 31) +
      (src31[3] << 31) +
      (src31[4] << 31) +
      (src31[5] << 31) +
      (src31[6] << 31) +
      (src31[7] << 31) +
      (src31[8] << 31) +
      (src31[9] << 31) +
      (src31[10] << 31) +
      (src31[11] << 31) +
      (src31[12] << 31) +
      (src31[13] << 31) +
      (src31[14] << 31) +
      (src31[15] << 31) +
      (src31[16] << 31) +
      (src31[17] << 31) +
      (src31[18] << 31) +
      (src31[19] << 31) +
      (src31[20] << 31) +
      (src31[21] << 31) +
      (src31[22] << 31) +
      (src31[23] << 31) +
      (src31[24] << 31) +
      (src31[25] << 31) +
      (src31[26] << 31) +
      (src31[27] << 31) +
      (src31[28] << 31) +
      (src31[29] << 31) +
      (src31[30] << 31) +
      (src31[31] << 31) +
      (src31[32] << 31) +
      (src31[33] << 31) +
      (src31[34] << 31) +
      (src31[35] << 31) +
      (src31[36] << 31) +
      (src31[37] << 31) +
      (src31[38] << 31) +
      (src31[39] << 31) +
      (src31[40] << 31) +
      (src31[41] << 31) +
      (src31[42] << 31) +
      (src31[43] << 31) +
      (src31[44] << 31) +
      (src31[45] << 31) +
      (src31[46] << 31) +
      (src31[47] << 31) +
      (src31[48] << 31) +
      (src31[49] << 31) +
      (src31[50] << 31) +
      (src31[51] << 31) +
      (src31[52] << 31) +
      (src31[53] << 31) +
      (src31[54] << 31) +
      (src31[55] << 31) +
      (src31[56] << 31) +
      (src31[57] << 31) +
      (src31[58] << 31) +
      (src31[59] << 31) +
      (src31[60] << 31) +
      (src31[61] << 31) +
      (src31[62] << 31) +
      (src31[63] << 31) +
      (src32[0] << 32) +
      (src32[1] << 32) +
      (src32[2] << 32) +
      (src32[3] << 32) +
      (src32[4] << 32) +
      (src32[5] << 32) +
      (src32[6] << 32) +
      (src32[7] << 32) +
      (src32[8] << 32) +
      (src32[9] << 32) +
      (src32[10] << 32) +
      (src32[11] << 32) +
      (src32[12] << 32) +
      (src32[13] << 32) +
      (src32[14] << 32) +
      (src32[15] << 32) +
      (src32[16] << 32) +
      (src32[17] << 32) +
      (src32[18] << 32) +
      (src32[19] << 32) +
      (src32[20] << 32) +
      (src32[21] << 32) +
      (src32[22] << 32) +
      (src32[23] << 32) +
      (src32[24] << 32) +
      (src32[25] << 32) +
      (src32[26] << 32) +
      (src32[27] << 32) +
      (src32[28] << 32) +
      (src32[29] << 32) +
      (src32[30] << 32) +
      (src32[31] << 32) +
      (src32[32] << 32) +
      (src32[33] << 32) +
      (src32[34] << 32) +
      (src32[35] << 32) +
      (src32[36] << 32) +
      (src32[37] << 32) +
      (src32[38] << 32) +
      (src32[39] << 32) +
      (src32[40] << 32) +
      (src32[41] << 32) +
      (src32[42] << 32) +
      (src32[43] << 32) +
      (src32[44] << 32) +
      (src32[45] << 32) +
      (src32[46] << 32) +
      (src32[47] << 32) +
      (src32[48] << 32) +
      (src32[49] << 32) +
      (src32[50] << 32) +
      (src32[51] << 32) +
      (src32[52] << 32) +
      (src32[53] << 32) +
      (src32[54] << 32) +
      (src32[55] << 32) +
      (src32[56] << 32) +
      (src32[57] << 32) +
      (src32[58] << 32) +
      (src32[59] << 32) +
      (src32[60] << 32) +
      (src32[61] << 32) +
      (src32[62] << 32) +
      (src32[63] << 32) +
      (src33[0] << 33) +
      (src33[1] << 33) +
      (src33[2] << 33) +
      (src33[3] << 33) +
      (src33[4] << 33) +
      (src33[5] << 33) +
      (src33[6] << 33) +
      (src33[7] << 33) +
      (src33[8] << 33) +
      (src33[9] << 33) +
      (src33[10] << 33) +
      (src33[11] << 33) +
      (src33[12] << 33) +
      (src33[13] << 33) +
      (src33[14] << 33) +
      (src33[15] << 33) +
      (src33[16] << 33) +
      (src33[17] << 33) +
      (src33[18] << 33) +
      (src33[19] << 33) +
      (src33[20] << 33) +
      (src33[21] << 33) +
      (src33[22] << 33) +
      (src33[23] << 33) +
      (src33[24] << 33) +
      (src33[25] << 33) +
      (src33[26] << 33) +
      (src33[27] << 33) +
      (src33[28] << 33) +
      (src33[29] << 33) +
      (src33[30] << 33) +
      (src33[31] << 33) +
      (src33[32] << 33) +
      (src33[33] << 33) +
      (src33[34] << 33) +
      (src33[35] << 33) +
      (src33[36] << 33) +
      (src33[37] << 33) +
      (src33[38] << 33) +
      (src33[39] << 33) +
      (src33[40] << 33) +
      (src33[41] << 33) +
      (src33[42] << 33) +
      (src33[43] << 33) +
      (src33[44] << 33) +
      (src33[45] << 33) +
      (src33[46] << 33) +
      (src33[47] << 33) +
      (src33[48] << 33) +
      (src33[49] << 33) +
      (src33[50] << 33) +
      (src33[51] << 33) +
      (src33[52] << 33) +
      (src33[53] << 33) +
      (src33[54] << 33) +
      (src33[55] << 33) +
      (src33[56] << 33) +
      (src33[57] << 33) +
      (src33[58] << 33) +
      (src33[59] << 33) +
      (src33[60] << 33) +
      (src33[61] << 33) +
      (src33[62] << 33) +
      (src33[63] << 33) +
      (src34[0] << 34) +
      (src34[1] << 34) +
      (src34[2] << 34) +
      (src34[3] << 34) +
      (src34[4] << 34) +
      (src34[5] << 34) +
      (src34[6] << 34) +
      (src34[7] << 34) +
      (src34[8] << 34) +
      (src34[9] << 34) +
      (src34[10] << 34) +
      (src34[11] << 34) +
      (src34[12] << 34) +
      (src34[13] << 34) +
      (src34[14] << 34) +
      (src34[15] << 34) +
      (src34[16] << 34) +
      (src34[17] << 34) +
      (src34[18] << 34) +
      (src34[19] << 34) +
      (src34[20] << 34) +
      (src34[21] << 34) +
      (src34[22] << 34) +
      (src34[23] << 34) +
      (src34[24] << 34) +
      (src34[25] << 34) +
      (src34[26] << 34) +
      (src34[27] << 34) +
      (src34[28] << 34) +
      (src34[29] << 34) +
      (src34[30] << 34) +
      (src34[31] << 34) +
      (src34[32] << 34) +
      (src34[33] << 34) +
      (src34[34] << 34) +
      (src34[35] << 34) +
      (src34[36] << 34) +
      (src34[37] << 34) +
      (src34[38] << 34) +
      (src34[39] << 34) +
      (src34[40] << 34) +
      (src34[41] << 34) +
      (src34[42] << 34) +
      (src34[43] << 34) +
      (src34[44] << 34) +
      (src34[45] << 34) +
      (src34[46] << 34) +
      (src34[47] << 34) +
      (src34[48] << 34) +
      (src34[49] << 34) +
      (src34[50] << 34) +
      (src34[51] << 34) +
      (src34[52] << 34) +
      (src34[53] << 34) +
      (src34[54] << 34) +
      (src34[55] << 34) +
      (src34[56] << 34) +
      (src34[57] << 34) +
      (src34[58] << 34) +
      (src34[59] << 34) +
      (src34[60] << 34) +
      (src34[61] << 34) +
      (src34[62] << 34) +
      (src34[63] << 34) +
      (src35[0] << 35) +
      (src35[1] << 35) +
      (src35[2] << 35) +
      (src35[3] << 35) +
      (src35[4] << 35) +
      (src35[5] << 35) +
      (src35[6] << 35) +
      (src35[7] << 35) +
      (src35[8] << 35) +
      (src35[9] << 35) +
      (src35[10] << 35) +
      (src35[11] << 35) +
      (src35[12] << 35) +
      (src35[13] << 35) +
      (src35[14] << 35) +
      (src35[15] << 35) +
      (src35[16] << 35) +
      (src35[17] << 35) +
      (src35[18] << 35) +
      (src35[19] << 35) +
      (src35[20] << 35) +
      (src35[21] << 35) +
      (src35[22] << 35) +
      (src35[23] << 35) +
      (src35[24] << 35) +
      (src35[25] << 35) +
      (src35[26] << 35) +
      (src35[27] << 35) +
      (src35[28] << 35) +
      (src35[29] << 35) +
      (src35[30] << 35) +
      (src35[31] << 35) +
      (src35[32] << 35) +
      (src35[33] << 35) +
      (src35[34] << 35) +
      (src35[35] << 35) +
      (src35[36] << 35) +
      (src35[37] << 35) +
      (src35[38] << 35) +
      (src35[39] << 35) +
      (src35[40] << 35) +
      (src35[41] << 35) +
      (src35[42] << 35) +
      (src35[43] << 35) +
      (src35[44] << 35) +
      (src35[45] << 35) +
      (src35[46] << 35) +
      (src35[47] << 35) +
      (src35[48] << 35) +
      (src35[49] << 35) +
      (src35[50] << 35) +
      (src35[51] << 35) +
      (src35[52] << 35) +
      (src35[53] << 35) +
      (src35[54] << 35) +
      (src35[55] << 35) +
      (src35[56] << 35) +
      (src35[57] << 35) +
      (src35[58] << 35) +
      (src35[59] << 35) +
      (src35[60] << 35) +
      (src35[61] << 35) +
      (src35[62] << 35) +
      (src35[63] << 35) +
      (src36[0] << 36) +
      (src36[1] << 36) +
      (src36[2] << 36) +
      (src36[3] << 36) +
      (src36[4] << 36) +
      (src36[5] << 36) +
      (src36[6] << 36) +
      (src36[7] << 36) +
      (src36[8] << 36) +
      (src36[9] << 36) +
      (src36[10] << 36) +
      (src36[11] << 36) +
      (src36[12] << 36) +
      (src36[13] << 36) +
      (src36[14] << 36) +
      (src36[15] << 36) +
      (src36[16] << 36) +
      (src36[17] << 36) +
      (src36[18] << 36) +
      (src36[19] << 36) +
      (src36[20] << 36) +
      (src36[21] << 36) +
      (src36[22] << 36) +
      (src36[23] << 36) +
      (src36[24] << 36) +
      (src36[25] << 36) +
      (src36[26] << 36) +
      (src36[27] << 36) +
      (src36[28] << 36) +
      (src36[29] << 36) +
      (src36[30] << 36) +
      (src36[31] << 36) +
      (src36[32] << 36) +
      (src36[33] << 36) +
      (src36[34] << 36) +
      (src36[35] << 36) +
      (src36[36] << 36) +
      (src36[37] << 36) +
      (src36[38] << 36) +
      (src36[39] << 36) +
      (src36[40] << 36) +
      (src36[41] << 36) +
      (src36[42] << 36) +
      (src36[43] << 36) +
      (src36[44] << 36) +
      (src36[45] << 36) +
      (src36[46] << 36) +
      (src36[47] << 36) +
      (src36[48] << 36) +
      (src36[49] << 36) +
      (src36[50] << 36) +
      (src36[51] << 36) +
      (src36[52] << 36) +
      (src36[53] << 36) +
      (src36[54] << 36) +
      (src36[55] << 36) +
      (src36[56] << 36) +
      (src36[57] << 36) +
      (src36[58] << 36) +
      (src36[59] << 36) +
      (src36[60] << 36) +
      (src36[61] << 36) +
      (src36[62] << 36) +
      (src36[63] << 36) +
      (src37[0] << 37) +
      (src37[1] << 37) +
      (src37[2] << 37) +
      (src37[3] << 37) +
      (src37[4] << 37) +
      (src37[5] << 37) +
      (src37[6] << 37) +
      (src37[7] << 37) +
      (src37[8] << 37) +
      (src37[9] << 37) +
      (src37[10] << 37) +
      (src37[11] << 37) +
      (src37[12] << 37) +
      (src37[13] << 37) +
      (src37[14] << 37) +
      (src37[15] << 37) +
      (src37[16] << 37) +
      (src37[17] << 37) +
      (src37[18] << 37) +
      (src37[19] << 37) +
      (src37[20] << 37) +
      (src37[21] << 37) +
      (src37[22] << 37) +
      (src37[23] << 37) +
      (src37[24] << 37) +
      (src37[25] << 37) +
      (src37[26] << 37) +
      (src37[27] << 37) +
      (src37[28] << 37) +
      (src37[29] << 37) +
      (src37[30] << 37) +
      (src37[31] << 37) +
      (src37[32] << 37) +
      (src37[33] << 37) +
      (src37[34] << 37) +
      (src37[35] << 37) +
      (src37[36] << 37) +
      (src37[37] << 37) +
      (src37[38] << 37) +
      (src37[39] << 37) +
      (src37[40] << 37) +
      (src37[41] << 37) +
      (src37[42] << 37) +
      (src37[43] << 37) +
      (src37[44] << 37) +
      (src37[45] << 37) +
      (src37[46] << 37) +
      (src37[47] << 37) +
      (src37[48] << 37) +
      (src37[49] << 37) +
      (src37[50] << 37) +
      (src37[51] << 37) +
      (src37[52] << 37) +
      (src37[53] << 37) +
      (src37[54] << 37) +
      (src37[55] << 37) +
      (src37[56] << 37) +
      (src37[57] << 37) +
      (src37[58] << 37) +
      (src37[59] << 37) +
      (src37[60] << 37) +
      (src37[61] << 37) +
      (src37[62] << 37) +
      (src37[63] << 37) +
      (src38[0] << 38) +
      (src38[1] << 38) +
      (src38[2] << 38) +
      (src38[3] << 38) +
      (src38[4] << 38) +
      (src38[5] << 38) +
      (src38[6] << 38) +
      (src38[7] << 38) +
      (src38[8] << 38) +
      (src38[9] << 38) +
      (src38[10] << 38) +
      (src38[11] << 38) +
      (src38[12] << 38) +
      (src38[13] << 38) +
      (src38[14] << 38) +
      (src38[15] << 38) +
      (src38[16] << 38) +
      (src38[17] << 38) +
      (src38[18] << 38) +
      (src38[19] << 38) +
      (src38[20] << 38) +
      (src38[21] << 38) +
      (src38[22] << 38) +
      (src38[23] << 38) +
      (src38[24] << 38) +
      (src38[25] << 38) +
      (src38[26] << 38) +
      (src38[27] << 38) +
      (src38[28] << 38) +
      (src38[29] << 38) +
      (src38[30] << 38) +
      (src38[31] << 38) +
      (src38[32] << 38) +
      (src38[33] << 38) +
      (src38[34] << 38) +
      (src38[35] << 38) +
      (src38[36] << 38) +
      (src38[37] << 38) +
      (src38[38] << 38) +
      (src38[39] << 38) +
      (src38[40] << 38) +
      (src38[41] << 38) +
      (src38[42] << 38) +
      (src38[43] << 38) +
      (src38[44] << 38) +
      (src38[45] << 38) +
      (src38[46] << 38) +
      (src38[47] << 38) +
      (src38[48] << 38) +
      (src38[49] << 38) +
      (src38[50] << 38) +
      (src38[51] << 38) +
      (src38[52] << 38) +
      (src38[53] << 38) +
      (src38[54] << 38) +
      (src38[55] << 38) +
      (src38[56] << 38) +
      (src38[57] << 38) +
      (src38[58] << 38) +
      (src38[59] << 38) +
      (src38[60] << 38) +
      (src38[61] << 38) +
      (src38[62] << 38) +
      (src38[63] << 38) +
      (src39[0] << 39) +
      (src39[1] << 39) +
      (src39[2] << 39) +
      (src39[3] << 39) +
      (src39[4] << 39) +
      (src39[5] << 39) +
      (src39[6] << 39) +
      (src39[7] << 39) +
      (src39[8] << 39) +
      (src39[9] << 39) +
      (src39[10] << 39) +
      (src39[11] << 39) +
      (src39[12] << 39) +
      (src39[13] << 39) +
      (src39[14] << 39) +
      (src39[15] << 39) +
      (src39[16] << 39) +
      (src39[17] << 39) +
      (src39[18] << 39) +
      (src39[19] << 39) +
      (src39[20] << 39) +
      (src39[21] << 39) +
      (src39[22] << 39) +
      (src39[23] << 39) +
      (src39[24] << 39) +
      (src39[25] << 39) +
      (src39[26] << 39) +
      (src39[27] << 39) +
      (src39[28] << 39) +
      (src39[29] << 39) +
      (src39[30] << 39) +
      (src39[31] << 39) +
      (src39[32] << 39) +
      (src39[33] << 39) +
      (src39[34] << 39) +
      (src39[35] << 39) +
      (src39[36] << 39) +
      (src39[37] << 39) +
      (src39[38] << 39) +
      (src39[39] << 39) +
      (src39[40] << 39) +
      (src39[41] << 39) +
      (src39[42] << 39) +
      (src39[43] << 39) +
      (src39[44] << 39) +
      (src39[45] << 39) +
      (src39[46] << 39) +
      (src39[47] << 39) +
      (src39[48] << 39) +
      (src39[49] << 39) +
      (src39[50] << 39) +
      (src39[51] << 39) +
      (src39[52] << 39) +
      (src39[53] << 39) +
      (src39[54] << 39) +
      (src39[55] << 39) +
      (src39[56] << 39) +
      (src39[57] << 39) +
      (src39[58] << 39) +
      (src39[59] << 39) +
      (src39[60] << 39) +
      (src39[61] << 39) +
      (src39[62] << 39) +
      (src39[63] << 39) +
      (src40[0] << 40) +
      (src40[1] << 40) +
      (src40[2] << 40) +
      (src40[3] << 40) +
      (src40[4] << 40) +
      (src40[5] << 40) +
      (src40[6] << 40) +
      (src40[7] << 40) +
      (src40[8] << 40) +
      (src40[9] << 40) +
      (src40[10] << 40) +
      (src40[11] << 40) +
      (src40[12] << 40) +
      (src40[13] << 40) +
      (src40[14] << 40) +
      (src40[15] << 40) +
      (src40[16] << 40) +
      (src40[17] << 40) +
      (src40[18] << 40) +
      (src40[19] << 40) +
      (src40[20] << 40) +
      (src40[21] << 40) +
      (src40[22] << 40) +
      (src40[23] << 40) +
      (src40[24] << 40) +
      (src40[25] << 40) +
      (src40[26] << 40) +
      (src40[27] << 40) +
      (src40[28] << 40) +
      (src40[29] << 40) +
      (src40[30] << 40) +
      (src40[31] << 40) +
      (src40[32] << 40) +
      (src40[33] << 40) +
      (src40[34] << 40) +
      (src40[35] << 40) +
      (src40[36] << 40) +
      (src40[37] << 40) +
      (src40[38] << 40) +
      (src40[39] << 40) +
      (src40[40] << 40) +
      (src40[41] << 40) +
      (src40[42] << 40) +
      (src40[43] << 40) +
      (src40[44] << 40) +
      (src40[45] << 40) +
      (src40[46] << 40) +
      (src40[47] << 40) +
      (src40[48] << 40) +
      (src40[49] << 40) +
      (src40[50] << 40) +
      (src40[51] << 40) +
      (src40[52] << 40) +
      (src40[53] << 40) +
      (src40[54] << 40) +
      (src40[55] << 40) +
      (src40[56] << 40) +
      (src40[57] << 40) +
      (src40[58] << 40) +
      (src40[59] << 40) +
      (src40[60] << 40) +
      (src40[61] << 40) +
      (src40[62] << 40) +
      (src40[63] << 40) +
      (src41[0] << 41) +
      (src41[1] << 41) +
      (src41[2] << 41) +
      (src41[3] << 41) +
      (src41[4] << 41) +
      (src41[5] << 41) +
      (src41[6] << 41) +
      (src41[7] << 41) +
      (src41[8] << 41) +
      (src41[9] << 41) +
      (src41[10] << 41) +
      (src41[11] << 41) +
      (src41[12] << 41) +
      (src41[13] << 41) +
      (src41[14] << 41) +
      (src41[15] << 41) +
      (src41[16] << 41) +
      (src41[17] << 41) +
      (src41[18] << 41) +
      (src41[19] << 41) +
      (src41[20] << 41) +
      (src41[21] << 41) +
      (src41[22] << 41) +
      (src41[23] << 41) +
      (src41[24] << 41) +
      (src41[25] << 41) +
      (src41[26] << 41) +
      (src41[27] << 41) +
      (src41[28] << 41) +
      (src41[29] << 41) +
      (src41[30] << 41) +
      (src41[31] << 41) +
      (src41[32] << 41) +
      (src41[33] << 41) +
      (src41[34] << 41) +
      (src41[35] << 41) +
      (src41[36] << 41) +
      (src41[37] << 41) +
      (src41[38] << 41) +
      (src41[39] << 41) +
      (src41[40] << 41) +
      (src41[41] << 41) +
      (src41[42] << 41) +
      (src41[43] << 41) +
      (src41[44] << 41) +
      (src41[45] << 41) +
      (src41[46] << 41) +
      (src41[47] << 41) +
      (src41[48] << 41) +
      (src41[49] << 41) +
      (src41[50] << 41) +
      (src41[51] << 41) +
      (src41[52] << 41) +
      (src41[53] << 41) +
      (src41[54] << 41) +
      (src41[55] << 41) +
      (src41[56] << 41) +
      (src41[57] << 41) +
      (src41[58] << 41) +
      (src41[59] << 41) +
      (src41[60] << 41) +
      (src41[61] << 41) +
      (src41[62] << 41) +
      (src41[63] << 41) +
      (src42[0] << 42) +
      (src42[1] << 42) +
      (src42[2] << 42) +
      (src42[3] << 42) +
      (src42[4] << 42) +
      (src42[5] << 42) +
      (src42[6] << 42) +
      (src42[7] << 42) +
      (src42[8] << 42) +
      (src42[9] << 42) +
      (src42[10] << 42) +
      (src42[11] << 42) +
      (src42[12] << 42) +
      (src42[13] << 42) +
      (src42[14] << 42) +
      (src42[15] << 42) +
      (src42[16] << 42) +
      (src42[17] << 42) +
      (src42[18] << 42) +
      (src42[19] << 42) +
      (src42[20] << 42) +
      (src42[21] << 42) +
      (src42[22] << 42) +
      (src42[23] << 42) +
      (src42[24] << 42) +
      (src42[25] << 42) +
      (src42[26] << 42) +
      (src42[27] << 42) +
      (src42[28] << 42) +
      (src42[29] << 42) +
      (src42[30] << 42) +
      (src42[31] << 42) +
      (src42[32] << 42) +
      (src42[33] << 42) +
      (src42[34] << 42) +
      (src42[35] << 42) +
      (src42[36] << 42) +
      (src42[37] << 42) +
      (src42[38] << 42) +
      (src42[39] << 42) +
      (src42[40] << 42) +
      (src42[41] << 42) +
      (src42[42] << 42) +
      (src42[43] << 42) +
      (src42[44] << 42) +
      (src42[45] << 42) +
      (src42[46] << 42) +
      (src42[47] << 42) +
      (src42[48] << 42) +
      (src42[49] << 42) +
      (src42[50] << 42) +
      (src42[51] << 42) +
      (src42[52] << 42) +
      (src42[53] << 42) +
      (src42[54] << 42) +
      (src42[55] << 42) +
      (src42[56] << 42) +
      (src42[57] << 42) +
      (src42[58] << 42) +
      (src42[59] << 42) +
      (src42[60] << 42) +
      (src42[61] << 42) +
      (src42[62] << 42) +
      (src42[63] << 42) +
      (src43[0] << 43) +
      (src43[1] << 43) +
      (src43[2] << 43) +
      (src43[3] << 43) +
      (src43[4] << 43) +
      (src43[5] << 43) +
      (src43[6] << 43) +
      (src43[7] << 43) +
      (src43[8] << 43) +
      (src43[9] << 43) +
      (src43[10] << 43) +
      (src43[11] << 43) +
      (src43[12] << 43) +
      (src43[13] << 43) +
      (src43[14] << 43) +
      (src43[15] << 43) +
      (src43[16] << 43) +
      (src43[17] << 43) +
      (src43[18] << 43) +
      (src43[19] << 43) +
      (src43[20] << 43) +
      (src43[21] << 43) +
      (src43[22] << 43) +
      (src43[23] << 43) +
      (src43[24] << 43) +
      (src43[25] << 43) +
      (src43[26] << 43) +
      (src43[27] << 43) +
      (src43[28] << 43) +
      (src43[29] << 43) +
      (src43[30] << 43) +
      (src43[31] << 43) +
      (src43[32] << 43) +
      (src43[33] << 43) +
      (src43[34] << 43) +
      (src43[35] << 43) +
      (src43[36] << 43) +
      (src43[37] << 43) +
      (src43[38] << 43) +
      (src43[39] << 43) +
      (src43[40] << 43) +
      (src43[41] << 43) +
      (src43[42] << 43) +
      (src43[43] << 43) +
      (src43[44] << 43) +
      (src43[45] << 43) +
      (src43[46] << 43) +
      (src43[47] << 43) +
      (src43[48] << 43) +
      (src43[49] << 43) +
      (src43[50] << 43) +
      (src43[51] << 43) +
      (src43[52] << 43) +
      (src43[53] << 43) +
      (src43[54] << 43) +
      (src43[55] << 43) +
      (src43[56] << 43) +
      (src43[57] << 43) +
      (src43[58] << 43) +
      (src43[59] << 43) +
      (src43[60] << 43) +
      (src43[61] << 43) +
      (src43[62] << 43) +
      (src43[63] << 43) +
      (src44[0] << 44) +
      (src44[1] << 44) +
      (src44[2] << 44) +
      (src44[3] << 44) +
      (src44[4] << 44) +
      (src44[5] << 44) +
      (src44[6] << 44) +
      (src44[7] << 44) +
      (src44[8] << 44) +
      (src44[9] << 44) +
      (src44[10] << 44) +
      (src44[11] << 44) +
      (src44[12] << 44) +
      (src44[13] << 44) +
      (src44[14] << 44) +
      (src44[15] << 44) +
      (src44[16] << 44) +
      (src44[17] << 44) +
      (src44[18] << 44) +
      (src44[19] << 44) +
      (src44[20] << 44) +
      (src44[21] << 44) +
      (src44[22] << 44) +
      (src44[23] << 44) +
      (src44[24] << 44) +
      (src44[25] << 44) +
      (src44[26] << 44) +
      (src44[27] << 44) +
      (src44[28] << 44) +
      (src44[29] << 44) +
      (src44[30] << 44) +
      (src44[31] << 44) +
      (src44[32] << 44) +
      (src44[33] << 44) +
      (src44[34] << 44) +
      (src44[35] << 44) +
      (src44[36] << 44) +
      (src44[37] << 44) +
      (src44[38] << 44) +
      (src44[39] << 44) +
      (src44[40] << 44) +
      (src44[41] << 44) +
      (src44[42] << 44) +
      (src44[43] << 44) +
      (src44[44] << 44) +
      (src44[45] << 44) +
      (src44[46] << 44) +
      (src44[47] << 44) +
      (src44[48] << 44) +
      (src44[49] << 44) +
      (src44[50] << 44) +
      (src44[51] << 44) +
      (src44[52] << 44) +
      (src44[53] << 44) +
      (src44[54] << 44) +
      (src44[55] << 44) +
      (src44[56] << 44) +
      (src44[57] << 44) +
      (src44[58] << 44) +
      (src44[59] << 44) +
      (src44[60] << 44) +
      (src44[61] << 44) +
      (src44[62] << 44) +
      (src44[63] << 44) +
      (src45[0] << 45) +
      (src45[1] << 45) +
      (src45[2] << 45) +
      (src45[3] << 45) +
      (src45[4] << 45) +
      (src45[5] << 45) +
      (src45[6] << 45) +
      (src45[7] << 45) +
      (src45[8] << 45) +
      (src45[9] << 45) +
      (src45[10] << 45) +
      (src45[11] << 45) +
      (src45[12] << 45) +
      (src45[13] << 45) +
      (src45[14] << 45) +
      (src45[15] << 45) +
      (src45[16] << 45) +
      (src45[17] << 45) +
      (src45[18] << 45) +
      (src45[19] << 45) +
      (src45[20] << 45) +
      (src45[21] << 45) +
      (src45[22] << 45) +
      (src45[23] << 45) +
      (src45[24] << 45) +
      (src45[25] << 45) +
      (src45[26] << 45) +
      (src45[27] << 45) +
      (src45[28] << 45) +
      (src45[29] << 45) +
      (src45[30] << 45) +
      (src45[31] << 45) +
      (src45[32] << 45) +
      (src45[33] << 45) +
      (src45[34] << 45) +
      (src45[35] << 45) +
      (src45[36] << 45) +
      (src45[37] << 45) +
      (src45[38] << 45) +
      (src45[39] << 45) +
      (src45[40] << 45) +
      (src45[41] << 45) +
      (src45[42] << 45) +
      (src45[43] << 45) +
      (src45[44] << 45) +
      (src45[45] << 45) +
      (src45[46] << 45) +
      (src45[47] << 45) +
      (src45[48] << 45) +
      (src45[49] << 45) +
      (src45[50] << 45) +
      (src45[51] << 45) +
      (src45[52] << 45) +
      (src45[53] << 45) +
      (src45[54] << 45) +
      (src45[55] << 45) +
      (src45[56] << 45) +
      (src45[57] << 45) +
      (src45[58] << 45) +
      (src45[59] << 45) +
      (src45[60] << 45) +
      (src45[61] << 45) +
      (src45[62] << 45) +
      (src45[63] << 45) +
      (src46[0] << 46) +
      (src46[1] << 46) +
      (src46[2] << 46) +
      (src46[3] << 46) +
      (src46[4] << 46) +
      (src46[5] << 46) +
      (src46[6] << 46) +
      (src46[7] << 46) +
      (src46[8] << 46) +
      (src46[9] << 46) +
      (src46[10] << 46) +
      (src46[11] << 46) +
      (src46[12] << 46) +
      (src46[13] << 46) +
      (src46[14] << 46) +
      (src46[15] << 46) +
      (src46[16] << 46) +
      (src46[17] << 46) +
      (src46[18] << 46) +
      (src46[19] << 46) +
      (src46[20] << 46) +
      (src46[21] << 46) +
      (src46[22] << 46) +
      (src46[23] << 46) +
      (src46[24] << 46) +
      (src46[25] << 46) +
      (src46[26] << 46) +
      (src46[27] << 46) +
      (src46[28] << 46) +
      (src46[29] << 46) +
      (src46[30] << 46) +
      (src46[31] << 46) +
      (src46[32] << 46) +
      (src46[33] << 46) +
      (src46[34] << 46) +
      (src46[35] << 46) +
      (src46[36] << 46) +
      (src46[37] << 46) +
      (src46[38] << 46) +
      (src46[39] << 46) +
      (src46[40] << 46) +
      (src46[41] << 46) +
      (src46[42] << 46) +
      (src46[43] << 46) +
      (src46[44] << 46) +
      (src46[45] << 46) +
      (src46[46] << 46) +
      (src46[47] << 46) +
      (src46[48] << 46) +
      (src46[49] << 46) +
      (src46[50] << 46) +
      (src46[51] << 46) +
      (src46[52] << 46) +
      (src46[53] << 46) +
      (src46[54] << 46) +
      (src46[55] << 46) +
      (src46[56] << 46) +
      (src46[57] << 46) +
      (src46[58] << 46) +
      (src46[59] << 46) +
      (src46[60] << 46) +
      (src46[61] << 46) +
      (src46[62] << 46) +
      (src46[63] << 46) +
      (src47[0] << 47) +
      (src47[1] << 47) +
      (src47[2] << 47) +
      (src47[3] << 47) +
      (src47[4] << 47) +
      (src47[5] << 47) +
      (src47[6] << 47) +
      (src47[7] << 47) +
      (src47[8] << 47) +
      (src47[9] << 47) +
      (src47[10] << 47) +
      (src47[11] << 47) +
      (src47[12] << 47) +
      (src47[13] << 47) +
      (src47[14] << 47) +
      (src47[15] << 47) +
      (src47[16] << 47) +
      (src47[17] << 47) +
      (src47[18] << 47) +
      (src47[19] << 47) +
      (src47[20] << 47) +
      (src47[21] << 47) +
      (src47[22] << 47) +
      (src47[23] << 47) +
      (src47[24] << 47) +
      (src47[25] << 47) +
      (src47[26] << 47) +
      (src47[27] << 47) +
      (src47[28] << 47) +
      (src47[29] << 47) +
      (src47[30] << 47) +
      (src47[31] << 47) +
      (src47[32] << 47) +
      (src47[33] << 47) +
      (src47[34] << 47) +
      (src47[35] << 47) +
      (src47[36] << 47) +
      (src47[37] << 47) +
      (src47[38] << 47) +
      (src47[39] << 47) +
      (src47[40] << 47) +
      (src47[41] << 47) +
      (src47[42] << 47) +
      (src47[43] << 47) +
      (src47[44] << 47) +
      (src47[45] << 47) +
      (src47[46] << 47) +
      (src47[47] << 47) +
      (src47[48] << 47) +
      (src47[49] << 47) +
      (src47[50] << 47) +
      (src47[51] << 47) +
      (src47[52] << 47) +
      (src47[53] << 47) +
      (src47[54] << 47) +
      (src47[55] << 47) +
      (src47[56] << 47) +
      (src47[57] << 47) +
      (src47[58] << 47) +
      (src47[59] << 47) +
      (src47[60] << 47) +
      (src47[61] << 47) +
      (src47[62] << 47) +
      (src47[63] << 47) +
      (src48[0] << 48) +
      (src48[1] << 48) +
      (src48[2] << 48) +
      (src48[3] << 48) +
      (src48[4] << 48) +
      (src48[5] << 48) +
      (src48[6] << 48) +
      (src48[7] << 48) +
      (src48[8] << 48) +
      (src48[9] << 48) +
      (src48[10] << 48) +
      (src48[11] << 48) +
      (src48[12] << 48) +
      (src48[13] << 48) +
      (src48[14] << 48) +
      (src48[15] << 48) +
      (src48[16] << 48) +
      (src48[17] << 48) +
      (src48[18] << 48) +
      (src48[19] << 48) +
      (src48[20] << 48) +
      (src48[21] << 48) +
      (src48[22] << 48) +
      (src48[23] << 48) +
      (src48[24] << 48) +
      (src48[25] << 48) +
      (src48[26] << 48) +
      (src48[27] << 48) +
      (src48[28] << 48) +
      (src48[29] << 48) +
      (src48[30] << 48) +
      (src48[31] << 48) +
      (src48[32] << 48) +
      (src48[33] << 48) +
      (src48[34] << 48) +
      (src48[35] << 48) +
      (src48[36] << 48) +
      (src48[37] << 48) +
      (src48[38] << 48) +
      (src48[39] << 48) +
      (src48[40] << 48) +
      (src48[41] << 48) +
      (src48[42] << 48) +
      (src48[43] << 48) +
      (src48[44] << 48) +
      (src48[45] << 48) +
      (src48[46] << 48) +
      (src48[47] << 48) +
      (src48[48] << 48) +
      (src48[49] << 48) +
      (src48[50] << 48) +
      (src48[51] << 48) +
      (src48[52] << 48) +
      (src48[53] << 48) +
      (src48[54] << 48) +
      (src48[55] << 48) +
      (src48[56] << 48) +
      (src48[57] << 48) +
      (src48[58] << 48) +
      (src48[59] << 48) +
      (src48[60] << 48) +
      (src48[61] << 48) +
      (src48[62] << 48) +
      (src48[63] << 48) +
      (src49[0] << 49) +
      (src49[1] << 49) +
      (src49[2] << 49) +
      (src49[3] << 49) +
      (src49[4] << 49) +
      (src49[5] << 49) +
      (src49[6] << 49) +
      (src49[7] << 49) +
      (src49[8] << 49) +
      (src49[9] << 49) +
      (src49[10] << 49) +
      (src49[11] << 49) +
      (src49[12] << 49) +
      (src49[13] << 49) +
      (src49[14] << 49) +
      (src49[15] << 49) +
      (src49[16] << 49) +
      (src49[17] << 49) +
      (src49[18] << 49) +
      (src49[19] << 49) +
      (src49[20] << 49) +
      (src49[21] << 49) +
      (src49[22] << 49) +
      (src49[23] << 49) +
      (src49[24] << 49) +
      (src49[25] << 49) +
      (src49[26] << 49) +
      (src49[27] << 49) +
      (src49[28] << 49) +
      (src49[29] << 49) +
      (src49[30] << 49) +
      (src49[31] << 49) +
      (src49[32] << 49) +
      (src49[33] << 49) +
      (src49[34] << 49) +
      (src49[35] << 49) +
      (src49[36] << 49) +
      (src49[37] << 49) +
      (src49[38] << 49) +
      (src49[39] << 49) +
      (src49[40] << 49) +
      (src49[41] << 49) +
      (src49[42] << 49) +
      (src49[43] << 49) +
      (src49[44] << 49) +
      (src49[45] << 49) +
      (src49[46] << 49) +
      (src49[47] << 49) +
      (src49[48] << 49) +
      (src49[49] << 49) +
      (src49[50] << 49) +
      (src49[51] << 49) +
      (src49[52] << 49) +
      (src49[53] << 49) +
      (src49[54] << 49) +
      (src49[55] << 49) +
      (src49[56] << 49) +
      (src49[57] << 49) +
      (src49[58] << 49) +
      (src49[59] << 49) +
      (src49[60] << 49) +
      (src49[61] << 49) +
      (src49[62] << 49) +
      (src49[63] << 49) +
      (src50[0] << 50) +
      (src50[1] << 50) +
      (src50[2] << 50) +
      (src50[3] << 50) +
      (src50[4] << 50) +
      (src50[5] << 50) +
      (src50[6] << 50) +
      (src50[7] << 50) +
      (src50[8] << 50) +
      (src50[9] << 50) +
      (src50[10] << 50) +
      (src50[11] << 50) +
      (src50[12] << 50) +
      (src50[13] << 50) +
      (src50[14] << 50) +
      (src50[15] << 50) +
      (src50[16] << 50) +
      (src50[17] << 50) +
      (src50[18] << 50) +
      (src50[19] << 50) +
      (src50[20] << 50) +
      (src50[21] << 50) +
      (src50[22] << 50) +
      (src50[23] << 50) +
      (src50[24] << 50) +
      (src50[25] << 50) +
      (src50[26] << 50) +
      (src50[27] << 50) +
      (src50[28] << 50) +
      (src50[29] << 50) +
      (src50[30] << 50) +
      (src50[31] << 50) +
      (src50[32] << 50) +
      (src50[33] << 50) +
      (src50[34] << 50) +
      (src50[35] << 50) +
      (src50[36] << 50) +
      (src50[37] << 50) +
      (src50[38] << 50) +
      (src50[39] << 50) +
      (src50[40] << 50) +
      (src50[41] << 50) +
      (src50[42] << 50) +
      (src50[43] << 50) +
      (src50[44] << 50) +
      (src50[45] << 50) +
      (src50[46] << 50) +
      (src50[47] << 50) +
      (src50[48] << 50) +
      (src50[49] << 50) +
      (src50[50] << 50) +
      (src50[51] << 50) +
      (src50[52] << 50) +
      (src50[53] << 50) +
      (src50[54] << 50) +
      (src50[55] << 50) +
      (src50[56] << 50) +
      (src50[57] << 50) +
      (src50[58] << 50) +
      (src50[59] << 50) +
      (src50[60] << 50) +
      (src50[61] << 50) +
      (src50[62] << 50) +
      (src50[63] << 50) +
      (src51[0] << 51) +
      (src51[1] << 51) +
      (src51[2] << 51) +
      (src51[3] << 51) +
      (src51[4] << 51) +
      (src51[5] << 51) +
      (src51[6] << 51) +
      (src51[7] << 51) +
      (src51[8] << 51) +
      (src51[9] << 51) +
      (src51[10] << 51) +
      (src51[11] << 51) +
      (src51[12] << 51) +
      (src51[13] << 51) +
      (src51[14] << 51) +
      (src51[15] << 51) +
      (src51[16] << 51) +
      (src51[17] << 51) +
      (src51[18] << 51) +
      (src51[19] << 51) +
      (src51[20] << 51) +
      (src51[21] << 51) +
      (src51[22] << 51) +
      (src51[23] << 51) +
      (src51[24] << 51) +
      (src51[25] << 51) +
      (src51[26] << 51) +
      (src51[27] << 51) +
      (src51[28] << 51) +
      (src51[29] << 51) +
      (src51[30] << 51) +
      (src51[31] << 51) +
      (src51[32] << 51) +
      (src51[33] << 51) +
      (src51[34] << 51) +
      (src51[35] << 51) +
      (src51[36] << 51) +
      (src51[37] << 51) +
      (src51[38] << 51) +
      (src51[39] << 51) +
      (src51[40] << 51) +
      (src51[41] << 51) +
      (src51[42] << 51) +
      (src51[43] << 51) +
      (src51[44] << 51) +
      (src51[45] << 51) +
      (src51[46] << 51) +
      (src51[47] << 51) +
      (src51[48] << 51) +
      (src51[49] << 51) +
      (src51[50] << 51) +
      (src51[51] << 51) +
      (src51[52] << 51) +
      (src51[53] << 51) +
      (src51[54] << 51) +
      (src51[55] << 51) +
      (src51[56] << 51) +
      (src51[57] << 51) +
      (src51[58] << 51) +
      (src51[59] << 51) +
      (src51[60] << 51) +
      (src51[61] << 51) +
      (src51[62] << 51) +
      (src51[63] << 51) +
      (src52[0] << 52) +
      (src52[1] << 52) +
      (src52[2] << 52) +
      (src52[3] << 52) +
      (src52[4] << 52) +
      (src52[5] << 52) +
      (src52[6] << 52) +
      (src52[7] << 52) +
      (src52[8] << 52) +
      (src52[9] << 52) +
      (src52[10] << 52) +
      (src52[11] << 52) +
      (src52[12] << 52) +
      (src52[13] << 52) +
      (src52[14] << 52) +
      (src52[15] << 52) +
      (src52[16] << 52) +
      (src52[17] << 52) +
      (src52[18] << 52) +
      (src52[19] << 52) +
      (src52[20] << 52) +
      (src52[21] << 52) +
      (src52[22] << 52) +
      (src52[23] << 52) +
      (src52[24] << 52) +
      (src52[25] << 52) +
      (src52[26] << 52) +
      (src52[27] << 52) +
      (src52[28] << 52) +
      (src52[29] << 52) +
      (src52[30] << 52) +
      (src52[31] << 52) +
      (src52[32] << 52) +
      (src52[33] << 52) +
      (src52[34] << 52) +
      (src52[35] << 52) +
      (src52[36] << 52) +
      (src52[37] << 52) +
      (src52[38] << 52) +
      (src52[39] << 52) +
      (src52[40] << 52) +
      (src52[41] << 52) +
      (src52[42] << 52) +
      (src52[43] << 52) +
      (src52[44] << 52) +
      (src52[45] << 52) +
      (src52[46] << 52) +
      (src52[47] << 52) +
      (src52[48] << 52) +
      (src52[49] << 52) +
      (src52[50] << 52) +
      (src52[51] << 52) +
      (src52[52] << 52) +
      (src52[53] << 52) +
      (src52[54] << 52) +
      (src52[55] << 52) +
      (src52[56] << 52) +
      (src52[57] << 52) +
      (src52[58] << 52) +
      (src52[59] << 52) +
      (src52[60] << 52) +
      (src52[61] << 52) +
      (src52[62] << 52) +
      (src52[63] << 52) +
      (src53[0] << 53) +
      (src53[1] << 53) +
      (src53[2] << 53) +
      (src53[3] << 53) +
      (src53[4] << 53) +
      (src53[5] << 53) +
      (src53[6] << 53) +
      (src53[7] << 53) +
      (src53[8] << 53) +
      (src53[9] << 53) +
      (src53[10] << 53) +
      (src53[11] << 53) +
      (src53[12] << 53) +
      (src53[13] << 53) +
      (src53[14] << 53) +
      (src53[15] << 53) +
      (src53[16] << 53) +
      (src53[17] << 53) +
      (src53[18] << 53) +
      (src53[19] << 53) +
      (src53[20] << 53) +
      (src53[21] << 53) +
      (src53[22] << 53) +
      (src53[23] << 53) +
      (src53[24] << 53) +
      (src53[25] << 53) +
      (src53[26] << 53) +
      (src53[27] << 53) +
      (src53[28] << 53) +
      (src53[29] << 53) +
      (src53[30] << 53) +
      (src53[31] << 53) +
      (src53[32] << 53) +
      (src53[33] << 53) +
      (src53[34] << 53) +
      (src53[35] << 53) +
      (src53[36] << 53) +
      (src53[37] << 53) +
      (src53[38] << 53) +
      (src53[39] << 53) +
      (src53[40] << 53) +
      (src53[41] << 53) +
      (src53[42] << 53) +
      (src53[43] << 53) +
      (src53[44] << 53) +
      (src53[45] << 53) +
      (src53[46] << 53) +
      (src53[47] << 53) +
      (src53[48] << 53) +
      (src53[49] << 53) +
      (src53[50] << 53) +
      (src53[51] << 53) +
      (src53[52] << 53) +
      (src53[53] << 53) +
      (src53[54] << 53) +
      (src53[55] << 53) +
      (src53[56] << 53) +
      (src53[57] << 53) +
      (src53[58] << 53) +
      (src53[59] << 53) +
      (src53[60] << 53) +
      (src53[61] << 53) +
      (src53[62] << 53) +
      (src53[63] << 53) +
      (src54[0] << 54) +
      (src54[1] << 54) +
      (src54[2] << 54) +
      (src54[3] << 54) +
      (src54[4] << 54) +
      (src54[5] << 54) +
      (src54[6] << 54) +
      (src54[7] << 54) +
      (src54[8] << 54) +
      (src54[9] << 54) +
      (src54[10] << 54) +
      (src54[11] << 54) +
      (src54[12] << 54) +
      (src54[13] << 54) +
      (src54[14] << 54) +
      (src54[15] << 54) +
      (src54[16] << 54) +
      (src54[17] << 54) +
      (src54[18] << 54) +
      (src54[19] << 54) +
      (src54[20] << 54) +
      (src54[21] << 54) +
      (src54[22] << 54) +
      (src54[23] << 54) +
      (src54[24] << 54) +
      (src54[25] << 54) +
      (src54[26] << 54) +
      (src54[27] << 54) +
      (src54[28] << 54) +
      (src54[29] << 54) +
      (src54[30] << 54) +
      (src54[31] << 54) +
      (src54[32] << 54) +
      (src54[33] << 54) +
      (src54[34] << 54) +
      (src54[35] << 54) +
      (src54[36] << 54) +
      (src54[37] << 54) +
      (src54[38] << 54) +
      (src54[39] << 54) +
      (src54[40] << 54) +
      (src54[41] << 54) +
      (src54[42] << 54) +
      (src54[43] << 54) +
      (src54[44] << 54) +
      (src54[45] << 54) +
      (src54[46] << 54) +
      (src54[47] << 54) +
      (src54[48] << 54) +
      (src54[49] << 54) +
      (src54[50] << 54) +
      (src54[51] << 54) +
      (src54[52] << 54) +
      (src54[53] << 54) +
      (src54[54] << 54) +
      (src54[55] << 54) +
      (src54[56] << 54) +
      (src54[57] << 54) +
      (src54[58] << 54) +
      (src54[59] << 54) +
      (src54[60] << 54) +
      (src54[61] << 54) +
      (src54[62] << 54) +
      (src54[63] << 54) +
      (src55[0] << 55) +
      (src55[1] << 55) +
      (src55[2] << 55) +
      (src55[3] << 55) +
      (src55[4] << 55) +
      (src55[5] << 55) +
      (src55[6] << 55) +
      (src55[7] << 55) +
      (src55[8] << 55) +
      (src55[9] << 55) +
      (src55[10] << 55) +
      (src55[11] << 55) +
      (src55[12] << 55) +
      (src55[13] << 55) +
      (src55[14] << 55) +
      (src55[15] << 55) +
      (src55[16] << 55) +
      (src55[17] << 55) +
      (src55[18] << 55) +
      (src55[19] << 55) +
      (src55[20] << 55) +
      (src55[21] << 55) +
      (src55[22] << 55) +
      (src55[23] << 55) +
      (src55[24] << 55) +
      (src55[25] << 55) +
      (src55[26] << 55) +
      (src55[27] << 55) +
      (src55[28] << 55) +
      (src55[29] << 55) +
      (src55[30] << 55) +
      (src55[31] << 55) +
      (src55[32] << 55) +
      (src55[33] << 55) +
      (src55[34] << 55) +
      (src55[35] << 55) +
      (src55[36] << 55) +
      (src55[37] << 55) +
      (src55[38] << 55) +
      (src55[39] << 55) +
      (src55[40] << 55) +
      (src55[41] << 55) +
      (src55[42] << 55) +
      (src55[43] << 55) +
      (src55[44] << 55) +
      (src55[45] << 55) +
      (src55[46] << 55) +
      (src55[47] << 55) +
      (src55[48] << 55) +
      (src55[49] << 55) +
      (src55[50] << 55) +
      (src55[51] << 55) +
      (src55[52] << 55) +
      (src55[53] << 55) +
      (src55[54] << 55) +
      (src55[55] << 55) +
      (src55[56] << 55) +
      (src55[57] << 55) +
      (src55[58] << 55) +
      (src55[59] << 55) +
      (src55[60] << 55) +
      (src55[61] << 55) +
      (src55[62] << 55) +
      (src55[63] << 55) +
      (src56[0] << 56) +
      (src56[1] << 56) +
      (src56[2] << 56) +
      (src56[3] << 56) +
      (src56[4] << 56) +
      (src56[5] << 56) +
      (src56[6] << 56) +
      (src56[7] << 56) +
      (src56[8] << 56) +
      (src56[9] << 56) +
      (src56[10] << 56) +
      (src56[11] << 56) +
      (src56[12] << 56) +
      (src56[13] << 56) +
      (src56[14] << 56) +
      (src56[15] << 56) +
      (src56[16] << 56) +
      (src56[17] << 56) +
      (src56[18] << 56) +
      (src56[19] << 56) +
      (src56[20] << 56) +
      (src56[21] << 56) +
      (src56[22] << 56) +
      (src56[23] << 56) +
      (src56[24] << 56) +
      (src56[25] << 56) +
      (src56[26] << 56) +
      (src56[27] << 56) +
      (src56[28] << 56) +
      (src56[29] << 56) +
      (src56[30] << 56) +
      (src56[31] << 56) +
      (src56[32] << 56) +
      (src56[33] << 56) +
      (src56[34] << 56) +
      (src56[35] << 56) +
      (src56[36] << 56) +
      (src56[37] << 56) +
      (src56[38] << 56) +
      (src56[39] << 56) +
      (src56[40] << 56) +
      (src56[41] << 56) +
      (src56[42] << 56) +
      (src56[43] << 56) +
      (src56[44] << 56) +
      (src56[45] << 56) +
      (src56[46] << 56) +
      (src56[47] << 56) +
      (src56[48] << 56) +
      (src56[49] << 56) +
      (src56[50] << 56) +
      (src56[51] << 56) +
      (src56[52] << 56) +
      (src56[53] << 56) +
      (src56[54] << 56) +
      (src56[55] << 56) +
      (src56[56] << 56) +
      (src56[57] << 56) +
      (src56[58] << 56) +
      (src56[59] << 56) +
      (src56[60] << 56) +
      (src56[61] << 56) +
      (src56[62] << 56) +
      (src56[63] << 56) +
      (src57[0] << 57) +
      (src57[1] << 57) +
      (src57[2] << 57) +
      (src57[3] << 57) +
      (src57[4] << 57) +
      (src57[5] << 57) +
      (src57[6] << 57) +
      (src57[7] << 57) +
      (src57[8] << 57) +
      (src57[9] << 57) +
      (src57[10] << 57) +
      (src57[11] << 57) +
      (src57[12] << 57) +
      (src57[13] << 57) +
      (src57[14] << 57) +
      (src57[15] << 57) +
      (src57[16] << 57) +
      (src57[17] << 57) +
      (src57[18] << 57) +
      (src57[19] << 57) +
      (src57[20] << 57) +
      (src57[21] << 57) +
      (src57[22] << 57) +
      (src57[23] << 57) +
      (src57[24] << 57) +
      (src57[25] << 57) +
      (src57[26] << 57) +
      (src57[27] << 57) +
      (src57[28] << 57) +
      (src57[29] << 57) +
      (src57[30] << 57) +
      (src57[31] << 57) +
      (src57[32] << 57) +
      (src57[33] << 57) +
      (src57[34] << 57) +
      (src57[35] << 57) +
      (src57[36] << 57) +
      (src57[37] << 57) +
      (src57[38] << 57) +
      (src57[39] << 57) +
      (src57[40] << 57) +
      (src57[41] << 57) +
      (src57[42] << 57) +
      (src57[43] << 57) +
      (src57[44] << 57) +
      (src57[45] << 57) +
      (src57[46] << 57) +
      (src57[47] << 57) +
      (src57[48] << 57) +
      (src57[49] << 57) +
      (src57[50] << 57) +
      (src57[51] << 57) +
      (src57[52] << 57) +
      (src57[53] << 57) +
      (src57[54] << 57) +
      (src57[55] << 57) +
      (src57[56] << 57) +
      (src57[57] << 57) +
      (src57[58] << 57) +
      (src57[59] << 57) +
      (src57[60] << 57) +
      (src57[61] << 57) +
      (src57[62] << 57) +
      (src57[63] << 57) +
      (src58[0] << 58) +
      (src58[1] << 58) +
      (src58[2] << 58) +
      (src58[3] << 58) +
      (src58[4] << 58) +
      (src58[5] << 58) +
      (src58[6] << 58) +
      (src58[7] << 58) +
      (src58[8] << 58) +
      (src58[9] << 58) +
      (src58[10] << 58) +
      (src58[11] << 58) +
      (src58[12] << 58) +
      (src58[13] << 58) +
      (src58[14] << 58) +
      (src58[15] << 58) +
      (src58[16] << 58) +
      (src58[17] << 58) +
      (src58[18] << 58) +
      (src58[19] << 58) +
      (src58[20] << 58) +
      (src58[21] << 58) +
      (src58[22] << 58) +
      (src58[23] << 58) +
      (src58[24] << 58) +
      (src58[25] << 58) +
      (src58[26] << 58) +
      (src58[27] << 58) +
      (src58[28] << 58) +
      (src58[29] << 58) +
      (src58[30] << 58) +
      (src58[31] << 58) +
      (src58[32] << 58) +
      (src58[33] << 58) +
      (src58[34] << 58) +
      (src58[35] << 58) +
      (src58[36] << 58) +
      (src58[37] << 58) +
      (src58[38] << 58) +
      (src58[39] << 58) +
      (src58[40] << 58) +
      (src58[41] << 58) +
      (src58[42] << 58) +
      (src58[43] << 58) +
      (src58[44] << 58) +
      (src58[45] << 58) +
      (src58[46] << 58) +
      (src58[47] << 58) +
      (src58[48] << 58) +
      (src58[49] << 58) +
      (src58[50] << 58) +
      (src58[51] << 58) +
      (src58[52] << 58) +
      (src58[53] << 58) +
      (src58[54] << 58) +
      (src58[55] << 58) +
      (src58[56] << 58) +
      (src58[57] << 58) +
      (src58[58] << 58) +
      (src58[59] << 58) +
      (src58[60] << 58) +
      (src58[61] << 58) +
      (src58[62] << 58) +
      (src58[63] << 58) +
      (src59[0] << 59) +
      (src59[1] << 59) +
      (src59[2] << 59) +
      (src59[3] << 59) +
      (src59[4] << 59) +
      (src59[5] << 59) +
      (src59[6] << 59) +
      (src59[7] << 59) +
      (src59[8] << 59) +
      (src59[9] << 59) +
      (src59[10] << 59) +
      (src59[11] << 59) +
      (src59[12] << 59) +
      (src59[13] << 59) +
      (src59[14] << 59) +
      (src59[15] << 59) +
      (src59[16] << 59) +
      (src59[17] << 59) +
      (src59[18] << 59) +
      (src59[19] << 59) +
      (src59[20] << 59) +
      (src59[21] << 59) +
      (src59[22] << 59) +
      (src59[23] << 59) +
      (src59[24] << 59) +
      (src59[25] << 59) +
      (src59[26] << 59) +
      (src59[27] << 59) +
      (src59[28] << 59) +
      (src59[29] << 59) +
      (src59[30] << 59) +
      (src59[31] << 59) +
      (src59[32] << 59) +
      (src59[33] << 59) +
      (src59[34] << 59) +
      (src59[35] << 59) +
      (src59[36] << 59) +
      (src59[37] << 59) +
      (src59[38] << 59) +
      (src59[39] << 59) +
      (src59[40] << 59) +
      (src59[41] << 59) +
      (src59[42] << 59) +
      (src59[43] << 59) +
      (src59[44] << 59) +
      (src59[45] << 59) +
      (src59[46] << 59) +
      (src59[47] << 59) +
      (src59[48] << 59) +
      (src59[49] << 59) +
      (src59[50] << 59) +
      (src59[51] << 59) +
      (src59[52] << 59) +
      (src59[53] << 59) +
      (src59[54] << 59) +
      (src59[55] << 59) +
      (src59[56] << 59) +
      (src59[57] << 59) +
      (src59[58] << 59) +
      (src59[59] << 59) +
      (src59[60] << 59) +
      (src59[61] << 59) +
      (src59[62] << 59) +
      (src59[63] << 59) +
      (src60[0] << 60) +
      (src60[1] << 60) +
      (src60[2] << 60) +
      (src60[3] << 60) +
      (src60[4] << 60) +
      (src60[5] << 60) +
      (src60[6] << 60) +
      (src60[7] << 60) +
      (src60[8] << 60) +
      (src60[9] << 60) +
      (src60[10] << 60) +
      (src60[11] << 60) +
      (src60[12] << 60) +
      (src60[13] << 60) +
      (src60[14] << 60) +
      (src60[15] << 60) +
      (src60[16] << 60) +
      (src60[17] << 60) +
      (src60[18] << 60) +
      (src60[19] << 60) +
      (src60[20] << 60) +
      (src60[21] << 60) +
      (src60[22] << 60) +
      (src60[23] << 60) +
      (src60[24] << 60) +
      (src60[25] << 60) +
      (src60[26] << 60) +
      (src60[27] << 60) +
      (src60[28] << 60) +
      (src60[29] << 60) +
      (src60[30] << 60) +
      (src60[31] << 60) +
      (src60[32] << 60) +
      (src60[33] << 60) +
      (src60[34] << 60) +
      (src60[35] << 60) +
      (src60[36] << 60) +
      (src60[37] << 60) +
      (src60[38] << 60) +
      (src60[39] << 60) +
      (src60[40] << 60) +
      (src60[41] << 60) +
      (src60[42] << 60) +
      (src60[43] << 60) +
      (src60[44] << 60) +
      (src60[45] << 60) +
      (src60[46] << 60) +
      (src60[47] << 60) +
      (src60[48] << 60) +
      (src60[49] << 60) +
      (src60[50] << 60) +
      (src60[51] << 60) +
      (src60[52] << 60) +
      (src60[53] << 60) +
      (src60[54] << 60) +
      (src60[55] << 60) +
      (src60[56] << 60) +
      (src60[57] << 60) +
      (src60[58] << 60) +
      (src60[59] << 60) +
      (src60[60] << 60) +
      (src60[61] << 60) +
      (src60[62] << 60) +
      (src60[63] << 60) +
      (src61[0] << 61) +
      (src61[1] << 61) +
      (src61[2] << 61) +
      (src61[3] << 61) +
      (src61[4] << 61) +
      (src61[5] << 61) +
      (src61[6] << 61) +
      (src61[7] << 61) +
      (src61[8] << 61) +
      (src61[9] << 61) +
      (src61[10] << 61) +
      (src61[11] << 61) +
      (src61[12] << 61) +
      (src61[13] << 61) +
      (src61[14] << 61) +
      (src61[15] << 61) +
      (src61[16] << 61) +
      (src61[17] << 61) +
      (src61[18] << 61) +
      (src61[19] << 61) +
      (src61[20] << 61) +
      (src61[21] << 61) +
      (src61[22] << 61) +
      (src61[23] << 61) +
      (src61[24] << 61) +
      (src61[25] << 61) +
      (src61[26] << 61) +
      (src61[27] << 61) +
      (src61[28] << 61) +
      (src61[29] << 61) +
      (src61[30] << 61) +
      (src61[31] << 61) +
      (src61[32] << 61) +
      (src61[33] << 61) +
      (src61[34] << 61) +
      (src61[35] << 61) +
      (src61[36] << 61) +
      (src61[37] << 61) +
      (src61[38] << 61) +
      (src61[39] << 61) +
      (src61[40] << 61) +
      (src61[41] << 61) +
      (src61[42] << 61) +
      (src61[43] << 61) +
      (src61[44] << 61) +
      (src61[45] << 61) +
      (src61[46] << 61) +
      (src61[47] << 61) +
      (src61[48] << 61) +
      (src61[49] << 61) +
      (src61[50] << 61) +
      (src61[51] << 61) +
      (src61[52] << 61) +
      (src61[53] << 61) +
      (src61[54] << 61) +
      (src61[55] << 61) +
      (src61[56] << 61) +
      (src61[57] << 61) +
      (src61[58] << 61) +
      (src61[59] << 61) +
      (src61[60] << 61) +
      (src61[61] << 61) +
      (src61[62] << 61) +
      (src61[63] << 61) +
      (src62[0] << 62) +
      (src62[1] << 62) +
      (src62[2] << 62) +
      (src62[3] << 62) +
      (src62[4] << 62) +
      (src62[5] << 62) +
      (src62[6] << 62) +
      (src62[7] << 62) +
      (src62[8] << 62) +
      (src62[9] << 62) +
      (src62[10] << 62) +
      (src62[11] << 62) +
      (src62[12] << 62) +
      (src62[13] << 62) +
      (src62[14] << 62) +
      (src62[15] << 62) +
      (src62[16] << 62) +
      (src62[17] << 62) +
      (src62[18] << 62) +
      (src62[19] << 62) +
      (src62[20] << 62) +
      (src62[21] << 62) +
      (src62[22] << 62) +
      (src62[23] << 62) +
      (src62[24] << 62) +
      (src62[25] << 62) +
      (src62[26] << 62) +
      (src62[27] << 62) +
      (src62[28] << 62) +
      (src62[29] << 62) +
      (src62[30] << 62) +
      (src62[31] << 62) +
      (src62[32] << 62) +
      (src62[33] << 62) +
      (src62[34] << 62) +
      (src62[35] << 62) +
      (src62[36] << 62) +
      (src62[37] << 62) +
      (src62[38] << 62) +
      (src62[39] << 62) +
      (src62[40] << 62) +
      (src62[41] << 62) +
      (src62[42] << 62) +
      (src62[43] << 62) +
      (src62[44] << 62) +
      (src62[45] << 62) +
      (src62[46] << 62) +
      (src62[47] << 62) +
      (src62[48] << 62) +
      (src62[49] << 62) +
      (src62[50] << 62) +
      (src62[51] << 62) +
      (src62[52] << 62) +
      (src62[53] << 62) +
      (src62[54] << 62) +
      (src62[55] << 62) +
      (src62[56] << 62) +
      (src62[57] << 62) +
      (src62[58] << 62) +
      (src62[59] << 62) +
      (src62[60] << 62) +
      (src62[61] << 62) +
      (src62[62] << 62) +
      (src62[63] << 62) +
      (src63[0] << 63) +
      (src63[1] << 63) +
      (src63[2] << 63) +
      (src63[3] << 63) +
      (src63[4] << 63) +
      (src63[5] << 63) +
      (src63[6] << 63) +
      (src63[7] << 63) +
      (src63[8] << 63) +
      (src63[9] << 63) +
      (src63[10] << 63) +
      (src63[11] << 63) +
      (src63[12] << 63) +
      (src63[13] << 63) +
      (src63[14] << 63) +
      (src63[15] << 63) +
      (src63[16] << 63) +
      (src63[17] << 63) +
      (src63[18] << 63) +
      (src63[19] << 63) +
      (src63[20] << 63) +
      (src63[21] << 63) +
      (src63[22] << 63) +
      (src63[23] << 63) +
      (src63[24] << 63) +
      (src63[25] << 63) +
      (src63[26] << 63) +
      (src63[27] << 63) +
      (src63[28] << 63) +
      (src63[29] << 63) +
      (src63[30] << 63) +
      (src63[31] << 63) +
      (src63[32] << 63) +
      (src63[33] << 63) +
      (src63[34] << 63) +
      (src63[35] << 63) +
      (src63[36] << 63) +
      (src63[37] << 63) +
      (src63[38] << 63) +
      (src63[39] << 63) +
      (src63[40] << 63) +
      (src63[41] << 63) +
      (src63[42] << 63) +
      (src63[43] << 63) +
      (src63[44] << 63) +
      (src63[45] << 63) +
      (src63[46] << 63) +
      (src63[47] << 63) +
      (src63[48] << 63) +
      (src63[49] << 63) +
      (src63[50] << 63) +
      (src63[51] << 63) +
      (src63[52] << 63) +
      (src63[53] << 63) +
      (src63[54] << 63) +
      (src63[55] << 63) +
      (src63[56] << 63) +
      (src63[57] << 63) +
      (src63[58] << 63) +
      (src63[59] << 63) +
      (src63[60] << 63) +
      (src63[61] << 63) +
      (src63[62] << 63) +
      (src63[63] << 63);
   assign dstsum =
      (dst00[0] << 0) +
      (dst00[1] << 0) +
      (dst01[0] << 1) +
      (dst02[0] << 2) +
      (dst02[1] << 2) +
      (dst03[0] << 3) +
      (dst03[1] << 3) +
      (dst04[0] << 4) +
      (dst04[1] << 4) +
      (dst05[0] << 5) +
      (dst05[1] << 5) +
      (dst06[0] << 6) +
      (dst06[1] << 6) +
      (dst07[0] << 7) +
      (dst07[1] << 7) +
      (dst08[0] << 8) +
      (dst09[0] << 9) +
      (dst09[1] << 9) +
      (dst10[0] << 10) +
      (dst10[1] << 10) +
      (dst11[0] << 11) +
      (dst11[1] << 11) +
      (dst12[0] << 12) +
      (dst12[1] << 12) +
      (dst13[0] << 13) +
      (dst13[1] << 13) +
      (dst14[0] << 14) +
      (dst14[1] << 14) +
      (dst15[0] << 15) +
      (dst15[1] << 15) +
      (dst16[0] << 16) +
      (dst16[1] << 16) +
      (dst17[0] << 17) +
      (dst17[1] << 17) +
      (dst18[0] << 18) +
      (dst18[1] << 18) +
      (dst19[0] << 19) +
      (dst19[1] << 19) +
      (dst20[0] << 20) +
      (dst21[0] << 21) +
      (dst21[1] << 21) +
      (dst22[0] << 22) +
      (dst22[1] << 22) +
      (dst23[0] << 23) +
      (dst23[1] << 23) +
      (dst24[0] << 24) +
      (dst24[1] << 24) +
      (dst25[0] << 25) +
      (dst25[1] << 25) +
      (dst26[0] << 26) +
      (dst26[1] << 26) +
      (dst27[0] << 27) +
      (dst27[1] << 27) +
      (dst28[0] << 28) +
      (dst28[1] << 28) +
      (dst29[0] << 29) +
      (dst29[1] << 29) +
      (dst30[0] << 30) +
      (dst30[1] << 30) +
      (dst31[0] << 31) +
      (dst32[0] << 32) +
      (dst32[1] << 32) +
      (dst33[0] << 33) +
      (dst33[1] << 33) +
      (dst34[0] << 34) +
      (dst35[0] << 35) +
      (dst35[1] << 35) +
      (dst36[0] << 36) +
      (dst36[1] << 36) +
      (dst37[0] << 37) +
      (dst37[1] << 37) +
      (dst38[0] << 38) +
      (dst38[1] << 38) +
      (dst39[0] << 39) +
      (dst39[1] << 39) +
      (dst40[0] << 40) +
      (dst40[1] << 40) +
      (dst41[0] << 41) +
      (dst41[1] << 41) +
      (dst42[0] << 42) +
      (dst42[1] << 42) +
      (dst43[0] << 43) +
      (dst43[1] << 43) +
      (dst44[0] << 44) +
      (dst44[1] << 44) +
      (dst45[0] << 45) +
      (dst45[1] << 45) +
      (dst46[0] << 46) +
      (dst47[0] << 47) +
      (dst47[1] << 47) +
      (dst48[0] << 48) +
      (dst48[1] << 48) +
      (dst49[0] << 49) +
      (dst49[1] << 49) +
      (dst50[0] << 50) +
      (dst50[1] << 50) +
      (dst51[0] << 51) +
      (dst51[1] << 51) +
      (dst52[0] << 52) +
      (dst52[1] << 52) +
      (dst53[0] << 53) +
      (dst53[1] << 53) +
      (dst54[0] << 54) +
      (dst54[1] << 54) +
      (dst55[0] << 55) +
      (dst55[1] << 55) +
      (dst56[0] << 56) +
      (dst56[1] << 56) +
      (dst57[0] << 57) +
      (dst57[1] << 57) +
      (dst58[0] << 58) +
      (dst59[0] << 59) +
      (dst59[1] << 59) +
      (dst60[0] << 60) +
      (dst60[1] << 60) +
      (dst61[0] << 61) +
      (dst61[1] << 61) +
      (dst62[0] << 62) +
      (dst62[1] << 62) +
      (dst63[0] << 63) +
      (dst63[1] << 63) +
      (dst64[0] << 64) +
      (dst65[0] << 65) +
      (dst65[1] << 65) +
      (dst66[0] << 66) +
      (dst66[1] << 66) +
      (dst67[0] << 67) +
      (dst67[1] << 67) +
      (dst68[0] << 68) +
      (dst68[1] << 68) +
      (dst69[0] << 69) +
      (dst69[1] << 69) +
      (dst70[0] << 70);
   compressor main_cmp(src00, src01, src02, src03, src04, src05, src06, src07, src08, src09, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, dst00, dst01, dst02, dst03, dst04, dst05, dst06, dst07, dst08, dst09, dst10, dst11, dst12, dst13, dst14, dst15, dst16, dst17, dst18, dst19, dst20, dst21, dst22, dst23, dst24, dst25, dst26, dst27, dst28, dst29, dst30, dst31, dst32, dst33, dst34, dst35, dst36, dst37, dst38, dst39, dst40, dst41, dst42, dst43, dst44, dst45, dst46, dst47, dst48, dst49, dst50, dst51, dst52, dst53, dst54, dst55, dst56, dst57, dst58, dst59, dst60, dst61, dst62, dst63, dst64, dst65, dst66, dst67, dst68, dst69, dst70);
   assign test = srcsum == dstsum;
   initial begin
      $monitor("src: 0x%x, dst: 0x%x, test: %b", srcsum, dstsum, test);
   end
   initial begin
      src00 <= 64'h0;
      src01 <= 64'h0;
      src02 <= 64'h0;
      src03 <= 64'h0;
      src04 <= 64'h0;
      src05 <= 64'h0;
      src06 <= 64'h0;
      src07 <= 64'h0;
      src08 <= 64'h0;
      src09 <= 64'h0;
      src10 <= 64'h0;
      src11 <= 64'h0;
      src12 <= 64'h0;
      src13 <= 64'h0;
      src14 <= 64'h0;
      src15 <= 64'h0;
      src16 <= 64'h0;
      src17 <= 64'h0;
      src18 <= 64'h0;
      src19 <= 64'h0;
      src20 <= 64'h0;
      src21 <= 64'h0;
      src22 <= 64'h0;
      src23 <= 64'h0;
      src24 <= 64'h0;
      src25 <= 64'h0;
      src26 <= 64'h0;
      src27 <= 64'h0;
      src28 <= 64'h0;
      src29 <= 64'h0;
      src30 <= 64'h0;
      src31 <= 64'h0;
      src32 <= 64'h0;
      src33 <= 64'h0;
      src34 <= 64'h0;
      src35 <= 64'h0;
      src36 <= 64'h0;
      src37 <= 64'h0;
      src38 <= 64'h0;
      src39 <= 64'h0;
      src40 <= 64'h0;
      src41 <= 64'h0;
      src42 <= 64'h0;
      src43 <= 64'h0;
      src44 <= 64'h0;
      src45 <= 64'h0;
      src46 <= 64'h0;
      src47 <= 64'h0;
      src48 <= 64'h0;
      src49 <= 64'h0;
      src50 <= 64'h0;
      src51 <= 64'h0;
      src52 <= 64'h0;
      src53 <= 64'h0;
      src54 <= 64'h0;
      src55 <= 64'h0;
      src56 <= 64'h0;
      src57 <= 64'h0;
      src58 <= 64'h0;
      src59 <= 64'h0;
      src60 <= 64'h0;
      src61 <= 64'h0;
      src62 <= 64'h0;
      src63 <= 64'h0;
      #1
      src00 <= 64'hffffffffffffffff;
      src01 <= 64'hffffffffffffffff;
      src02 <= 64'hffffffffffffffff;
      src03 <= 64'hffffffffffffffff;
      src04 <= 64'hffffffffffffffff;
      src05 <= 64'hffffffffffffffff;
      src06 <= 64'hffffffffffffffff;
      src07 <= 64'hffffffffffffffff;
      src08 <= 64'hffffffffffffffff;
      src09 <= 64'hffffffffffffffff;
      src10 <= 64'hffffffffffffffff;
      src11 <= 64'hffffffffffffffff;
      src12 <= 64'hffffffffffffffff;
      src13 <= 64'hffffffffffffffff;
      src14 <= 64'hffffffffffffffff;
      src15 <= 64'hffffffffffffffff;
      src16 <= 64'hffffffffffffffff;
      src17 <= 64'hffffffffffffffff;
      src18 <= 64'hffffffffffffffff;
      src19 <= 64'hffffffffffffffff;
      src20 <= 64'hffffffffffffffff;
      src21 <= 64'hffffffffffffffff;
      src22 <= 64'hffffffffffffffff;
      src23 <= 64'hffffffffffffffff;
      src24 <= 64'hffffffffffffffff;
      src25 <= 64'hffffffffffffffff;
      src26 <= 64'hffffffffffffffff;
      src27 <= 64'hffffffffffffffff;
      src28 <= 64'hffffffffffffffff;
      src29 <= 64'hffffffffffffffff;
      src30 <= 64'hffffffffffffffff;
      src31 <= 64'hffffffffffffffff;
      src32 <= 64'hffffffffffffffff;
      src33 <= 64'hffffffffffffffff;
      src34 <= 64'hffffffffffffffff;
      src35 <= 64'hffffffffffffffff;
      src36 <= 64'hffffffffffffffff;
      src37 <= 64'hffffffffffffffff;
      src38 <= 64'hffffffffffffffff;
      src39 <= 64'hffffffffffffffff;
      src40 <= 64'hffffffffffffffff;
      src41 <= 64'hffffffffffffffff;
      src42 <= 64'hffffffffffffffff;
      src43 <= 64'hffffffffffffffff;
      src44 <= 64'hffffffffffffffff;
      src45 <= 64'hffffffffffffffff;
      src46 <= 64'hffffffffffffffff;
      src47 <= 64'hffffffffffffffff;
      src48 <= 64'hffffffffffffffff;
      src49 <= 64'hffffffffffffffff;
      src50 <= 64'hffffffffffffffff;
      src51 <= 64'hffffffffffffffff;
      src52 <= 64'hffffffffffffffff;
      src53 <= 64'hffffffffffffffff;
      src54 <= 64'hffffffffffffffff;
      src55 <= 64'hffffffffffffffff;
      src56 <= 64'hffffffffffffffff;
      src57 <= 64'hffffffffffffffff;
      src58 <= 64'hffffffffffffffff;
      src59 <= 64'hffffffffffffffff;
      src60 <= 64'hffffffffffffffff;
      src61 <= 64'hffffffffffffffff;
      src62 <= 64'hffffffffffffffff;
      src63 <= 64'hffffffffffffffff;
      #1
      src00 <= 64'h6baa9455e3e70682;
      src01 <= 64'hd4713d60c8a70639;
      src02 <= 64'h7a024204f7c1bd87;
      src03 <= 64'h8133287637ebdcd9;
      src04 <= 64'h4f65d4d9259f4329;
      src05 <= 64'haf19922ad9b8a714;
      src06 <= 64'h8f4ff31e78de5857;
      src07 <= 64'h6f25e2a25a921187;
      src08 <= 64'h42af9fc385776e9a;
      src09 <= 64'h3983ca8ea7e9d49;
      src10 <= 64'hd71037d1b83e90ec;
      src11 <= 64'ha0116be5ab0c1681;
      src12 <= 64'h55485822de1b372a;
      src13 <= 64'h101fbcccded733e8;
      src14 <= 64'h9148624feac1c14f;
      src15 <= 64'h1759edc372ae2244;
      src16 <= 64'h1beb37117d41e602;
      src17 <= 64'h8c25166a1ff39849;
      src18 <= 64'h71eacd0549a3e80e;
      src19 <= 64'hcc45782198a6416d;
      src20 <= 64'h935ddd725129fb7c;
      src21 <= 64'h2f1205544a5308cc;
      src22 <= 64'h2fcd81b5d24bace4;
      src23 <= 64'h79fdef7c42930b33;
      src24 <= 64'he07405eb215663ab;
      src25 <= 64'h864a7a50b48d73f1;
      src26 <= 64'hcfc6e62585940927;
      src27 <= 64'h73581a8146743741;
      src28 <= 64'h5b7c709acb175a5a;
      src29 <= 64'h9cdf5a865306f3f5;
      src30 <= 64'hd857010255d44936;
      src31 <= 64'h552116dd2ba4b180;
      src32 <= 64'hfebd845d0dfae43;
      src33 <= 64'h38018b47b29a8b06;
      src34 <= 64'hae3b16ec9a27d858;
      src35 <= 64'h1ea45cd69371a71f;
      src36 <= 64'h1db53334fb0323a1;
      src37 <= 64'h589f8779b025244;
      src38 <= 64'hf87f43fdf6062541;
      src39 <= 64'h1fb797fab7d6467b;
      src40 <= 64'h8b53031d05d51433;
      src41 <= 64'h11ebcd49428a1c22;
      src42 <= 64'ha59cec98126cbc8f;
      src43 <= 64'h6fa231e959acdd98;
      src44 <= 64'h80ee526e0fa07a3f;
      src45 <= 64'h98b33c6e0a14b90a;
      src46 <= 64'hfcfcfa81b306d700;
      src47 <= 64'h429817c53308fb2e;
      src48 <= 64'hbb4a06cbe786ab37;
      src49 <= 64'h361524c2cc0f859;
      src50 <= 64'h403d1f83a859890c;
      src51 <= 64'hb0d9c2aa8f837ef7;
      src52 <= 64'hbdd7d19b753c7c99;
      src53 <= 64'hbd30291a55fea08e;
      src54 <= 64'h47e7f5938b5885ca;
      src55 <= 64'hac642b4c49b25ded;
      src56 <= 64'hb732d46f21e15094;
      src57 <= 64'hbf9cc545635518f7;
      src58 <= 64'ha69cfb85d432f8db;
      src59 <= 64'h983631890063e42f;
      src60 <= 64'h559b5975b2d650af;
      src61 <= 64'h6a1689addfe1b307;
      src62 <= 64'hb5816b74a985ab61;
      src63 <= 64'h720299e32a69acc7;
      #1
      src00 <= 64'hb3969057425cb200;
      src01 <= 64'hc167733f9a9e4310;
      src02 <= 64'h9f6048fe245a460;
      src03 <= 64'h6a46721acffa6cdd;
      src04 <= 64'hfa83ada4a2121ac5;
      src05 <= 64'hb9bdee2dd663049d;
      src06 <= 64'h3c54c71fca05536;
      src07 <= 64'hadb328cbf3158c0c;
      src08 <= 64'hde59f550f0fc2b;
      src09 <= 64'h30c1fb6a19086515;
      src10 <= 64'ha636425c9bbd750d;
      src11 <= 64'h4d6b234fdfa7c6ed;
      src12 <= 64'hfa7ff8bfb044284a;
      src13 <= 64'h597aab614d30dbc;
      src14 <= 64'h58d87776a51ad4f3;
      src15 <= 64'h27896389df3277fd;
      src16 <= 64'h4c14982d9ead926;
      src17 <= 64'h8ef066d44279b14d;
      src18 <= 64'he7180322a4e695c9;
      src19 <= 64'h6f790959a3e04b3b;
      src20 <= 64'h89b5b368df14c612;
      src21 <= 64'h247145f4a814d53;
      src22 <= 64'h4578bab326a97465;
      src23 <= 64'hca24be4d56672017;
      src24 <= 64'h17fd3736b7ef941c;
      src25 <= 64'h9edb95f2c787ddfb;
      src26 <= 64'h4505f4f60a8c46c7;
      src27 <= 64'h5c6460364a1eb1b7;
      src28 <= 64'h8c69778ffd42f697;
      src29 <= 64'h1d69d9fc4b1cb8bd;
      src30 <= 64'h4ed135530c5a876f;
      src31 <= 64'h4d7bd307122411e6;
      src32 <= 64'h5419eefcd5e73e3f;
      src33 <= 64'h1bd094486a2b3200;
      src34 <= 64'he89dc8158f928dc5;
      src35 <= 64'h1fd3c01757f98d1e;
      src36 <= 64'hb318ad4c1db2b452;
      src37 <= 64'h9aedbd06d316b4a;
      src38 <= 64'ha38d8afcfdd2ed7a;
      src39 <= 64'hceca2ee310da8a95;
      src40 <= 64'hbff773ce32b2c492;
      src41 <= 64'h628308690fa7ee05;
      src42 <= 64'h4a31b24384dd6da6;
      src43 <= 64'h6c4c3935379deda1;
      src44 <= 64'h2aa50f4ec6f00933;
      src45 <= 64'h5bc7fdeb31234efe;
      src46 <= 64'hb3b68b57da54f267;
      src47 <= 64'h869bdbd2e72bb5b7;
      src48 <= 64'had4ab155c09fcd8f;
      src49 <= 64'h7f411fed1e70e799;
      src50 <= 64'h1ac902ee25777cf0;
      src51 <= 64'h60c6b3ed755a3ac1;
      src52 <= 64'hd3b564b08be04c3e;
      src53 <= 64'h7ce71b48fba52e59;
      src54 <= 64'he345ac72eac39204;
      src55 <= 64'hee6a8e2f9c19ed34;
      src56 <= 64'hd17034ce51797350;
      src57 <= 64'h866d7002091472ad;
      src58 <= 64'h953c178e61067a8c;
      src59 <= 64'ha1727f7ea5f24b6;
      src60 <= 64'h21681081399f8a8f;
      src61 <= 64'h72d6bc20d80d6a1c;
      src62 <= 64'hf7f60e7f75f2bc20;
      src63 <= 64'h809f292387a1798f;
      #1
      src00 <= 64'hbf391fbb138c3460;
      src01 <= 64'hc12ea9b8e7e13ed8;
      src02 <= 64'hf8e45086ca819c6f;
      src03 <= 64'h961d8dcf9b8086da;
      src04 <= 64'hbda17da2000fc63d;
      src05 <= 64'h552ae5ca4124405b;
      src06 <= 64'hdc2151e17e56ac3d;
      src07 <= 64'hd334886ff164f9d8;
      src08 <= 64'h68777babc5c14262;
      src09 <= 64'h6238d0a0cf5e9ea3;
      src10 <= 64'h3d2bf042209818d1;
      src11 <= 64'hd476fe38babd4745;
      src12 <= 64'hf11ddff70e370526;
      src13 <= 64'h6af944e07b38785b;
      src14 <= 64'hb799ae8e9a1a7d6f;
      src15 <= 64'hb2ddc481ac6d5df8;
      src16 <= 64'hfc98c279cf6f111c;
      src17 <= 64'h62fda854775e0ec3;
      src18 <= 64'h19faa06e0c0a5967;
      src19 <= 64'h26c00984c734bb05;
      src20 <= 64'ha145789921f8c156;
      src21 <= 64'h58bf3b9ea6245b59;
      src22 <= 64'h7d859725c707aef9;
      src23 <= 64'hef151673a1df3da7;
      src24 <= 64'hcca1a034633cbf79;
      src25 <= 64'h71cff814645bd776;
      src26 <= 64'h30c32323c1b199c4;
      src27 <= 64'hf4dd05d51349747a;
      src28 <= 64'hef2d9a38e6e4b8df;
      src29 <= 64'h374a6cc9e0397e67;
      src30 <= 64'hf20b575d4e28e674;
      src31 <= 64'hef8d9ff015831fee;
      src32 <= 64'h101bb5fa6a677623;
      src33 <= 64'hc618fc1e6a480542;
      src34 <= 64'hf45da406bbf9bb01;
      src35 <= 64'h725c2675ca9571e4;
      src36 <= 64'h6ac1ca75afb918c8;
      src37 <= 64'h141b1a1b40a978bf;
      src38 <= 64'h1f12a0e912011caa;
      src39 <= 64'h78548d7b1182d23;
      src40 <= 64'h2d8b5b41590e83da;
      src41 <= 64'hf96d4403d48c93f3;
      src42 <= 64'h5da53b38d1aa6c5e;
      src43 <= 64'he4b8298798ba0f0e;
      src44 <= 64'hd3d1af353e0c86;
      src45 <= 64'he6a1a40bf031f4b9;
      src46 <= 64'h1d6d903bf7b68ae;
      src47 <= 64'hb080e0035e7f503c;
      src48 <= 64'h9ad7558feecb325b;
      src49 <= 64'h2452bc39dbf2eed1;
      src50 <= 64'h1cc5a8a0743c7e9d;
      src51 <= 64'h215203c7421aa15e;
      src52 <= 64'h35475c5ef76dce6e;
      src53 <= 64'h53b53b92a2cb5f38;
      src54 <= 64'hfe3216bd97d01e70;
      src55 <= 64'h280a07ee4ec985ff;
      src56 <= 64'hcdec85da200f7753;
      src57 <= 64'h8222134550de4292;
      src58 <= 64'hc13e66af3c9590d3;
      src59 <= 64'h5f59aa2c4a82e06a;
      src60 <= 64'h99e8c82821da132c;
      src61 <= 64'h21cc14b312bdf75f;
      src62 <= 64'h8cffbbb14ca49aaf;
      src63 <= 64'hed28508dbdaa3bfa;
      #1
      src00 <= 64'h6c148fc69750ca7e;
      src01 <= 64'h5ac4b6c7a31034dd;
      src02 <= 64'hecfb95b877a2133;
      src03 <= 64'h2284fd9689bba65;
      src04 <= 64'h70f8dd9952177eb7;
      src05 <= 64'hcbe88a3f2f7a304f;
      src06 <= 64'hb02de52c9b050db2;
      src07 <= 64'hb3dd77e1cbb02fe9;
      src08 <= 64'h66163e5beda2fc4c;
      src09 <= 64'h6bf4d047c4841a8d;
      src10 <= 64'h247f4d9785fa2d5c;
      src11 <= 64'h4b7350d13421beaf;
      src12 <= 64'hb2f11ef9d4864482;
      src13 <= 64'h764657ca9e65736c;
      src14 <= 64'h4c6e6fbb37fef6b5;
      src15 <= 64'h78aff58ec058a332;
      src16 <= 64'h67c21355c3121af6;
      src17 <= 64'hfbe86a8ea1cf0d1d;
      src18 <= 64'ha614be3ab2212c9;
      src19 <= 64'h71d04b0f656fa7e6;
      src20 <= 64'h40aaec7abf1df687;
      src21 <= 64'he8a56f31ac2c10d0;
      src22 <= 64'h15d38ca9986cc8d5;
      src23 <= 64'hcad00273120961ea;
      src24 <= 64'h889c8ae24e3c0f2d;
      src25 <= 64'h29deb984c31277fd;
      src26 <= 64'hdc66a27b6a325333;
      src27 <= 64'h8513d91e48622a67;
      src28 <= 64'h88083ebc35d4cd35;
      src29 <= 64'h4ad12b4c47534952;
      src30 <= 64'h2835bcdb2347b24f;
      src31 <= 64'h1eda4209b270af55;
      src32 <= 64'h974fdedc66b62087;
      src33 <= 64'hbe0a5a5679009c61;
      src34 <= 64'h7a0a02ba37cf8025;
      src35 <= 64'h8066b49bb1d792a0;
      src36 <= 64'h71a8c9c60f6ab75b;
      src37 <= 64'hbec60ffe248f4a25;
      src38 <= 64'h68a3c383739076a;
      src39 <= 64'hfa999f9b86de3365;
      src40 <= 64'hddfae808afd86432;
      src41 <= 64'hab4414aeecb3d561;
      src42 <= 64'h5c7cbc6201a4f7a1;
      src43 <= 64'h9ef1c8461dbc24fd;
      src44 <= 64'hb31e9be8a3ef802e;
      src45 <= 64'he695f8baba2338fe;
      src46 <= 64'h30f2c48549b564fb;
      src47 <= 64'h62565a955487b5c3;
      src48 <= 64'haffe2554e5aef699;
      src49 <= 64'h2114c2d650ea1324;
      src50 <= 64'h2fd3b9f2e90f79f8;
      src51 <= 64'hcbab5b51385c5fdc;
      src52 <= 64'hf0a61c5e707421d4;
      src53 <= 64'hb5c25d429626d8c4;
      src54 <= 64'h636abf8ce7e3f52c;
      src55 <= 64'ha217cf253be95767;
      src56 <= 64'h2fcf3b87defa7864;
      src57 <= 64'h2c623ac3ad7027cf;
      src58 <= 64'hc061c99b831a352a;
      src59 <= 64'h6953a1155a62ddc4;
      src60 <= 64'h94b9cdb56e3c18c9;
      src61 <= 64'h3725bd0c79c45c38;
      src62 <= 64'hacfeba4441030ae;
      src63 <= 64'h29b108230d742256;
      #1
      src00 <= 64'h23f1b67e01d34690;
      src01 <= 64'h7425f4e93891aef5;
      src02 <= 64'h9bbac83856e9b78d;
      src03 <= 64'he2014a459b3a0c89;
      src04 <= 64'h51abf5e5cb775e24;
      src05 <= 64'h4168705a533c9a31;
      src06 <= 64'hb5aafef85a1282a;
      src07 <= 64'h14827a895e6364c6;
      src08 <= 64'h864696c1deb4e6c4;
      src09 <= 64'hd658b1b33012ae1c;
      src10 <= 64'h4d236555bc5074ac;
      src11 <= 64'hdc2897c684539813;
      src12 <= 64'h7b69e69041300879;
      src13 <= 64'hb6651d6edf39ccaa;
      src14 <= 64'h1284b9d78d4e2753;
      src15 <= 64'h75e417dd7e5b637d;
      src16 <= 64'h15eae9d21e3d59d0;
      src17 <= 64'h275f275cc3f3f74d;
      src18 <= 64'heb52ee01e25e6512;
      src19 <= 64'h9cdd9f6c70cdc4a8;
      src20 <= 64'h3fee2fc72e2dffdf;
      src21 <= 64'hc9fe60368a83efc8;
      src22 <= 64'h45c596d442d01ba3;
      src23 <= 64'hb63f83c6c89309e9;
      src24 <= 64'hbb9e5a022c2df3c2;
      src25 <= 64'h37d316a43fafa217;
      src26 <= 64'h83e9973b89181ba3;
      src27 <= 64'hcbdc014dbedb42e;
      src28 <= 64'ha52ba0ce627b585f;
      src29 <= 64'h5be12d09908e0372;
      src30 <= 64'ha91da2cd8bf06f64;
      src31 <= 64'h3d798f0be6cd3595;
      src32 <= 64'h3bcd6aec53ca8c05;
      src33 <= 64'h7af2f402a0e624f1;
      src34 <= 64'h2bdfb7279501e917;
      src35 <= 64'h53f04099813dd49a;
      src36 <= 64'ha283453695decd6e;
      src37 <= 64'hd0f0c75d21d32e24;
      src38 <= 64'h62759469c28d2ad5;
      src39 <= 64'h974d9d499bc69882;
      src40 <= 64'h5bce228b989bb030;
      src41 <= 64'h4f06ea1874a26444;
      src42 <= 64'hbcc4616df40d2a37;
      src43 <= 64'h142a6c95d9082a42;
      src44 <= 64'h9ab3cc27232f8c5b;
      src45 <= 64'hc90ded295100f186;
      src46 <= 64'hf19b43da6253dfe3;
      src47 <= 64'h9cd3bdf356af737;
      src48 <= 64'ha867a0f0a8e6a772;
      src49 <= 64'h4e0e15d3298e9a79;
      src50 <= 64'h5a79b46a26b61b06;
      src51 <= 64'ha0b976c27db931ce;
      src52 <= 64'h3dd0c8660649def5;
      src53 <= 64'h53a081a6a7647989;
      src54 <= 64'hff9d318d22a3a62;
      src55 <= 64'ha9fa4ea6f8db1a4d;
      src56 <= 64'h72ef7dce376e22a6;
      src57 <= 64'h5ba830dc245db6ca;
      src58 <= 64'ha629d3322d4ba5a4;
      src59 <= 64'h689c0559bf4fa4a3;
      src60 <= 64'hb476998dafc8128a;
      src61 <= 64'h1f626a97ebe7ef91;
      src62 <= 64'h63eaa07ff436498e;
      src63 <= 64'h8024532000cbd313;
      #1
      src00 <= 64'h25ee54abb3191702;
      src01 <= 64'hd216ad53d4088ff7;
      src02 <= 64'hf22a4fc63f2de8a8;
      src03 <= 64'hb7c144fb2b16ad04;
      src04 <= 64'h40a210150a40a379;
      src05 <= 64'he3b4df81eeb3462c;
      src06 <= 64'h16f14aad7f107645;
      src07 <= 64'habf0f4bd4af0a6fe;
      src08 <= 64'h679b29e8c0c32da9;
      src09 <= 64'hcda6a326451437d6;
      src10 <= 64'h6480fdc0f1c58f44;
      src11 <= 64'h8cea309b49c94aa5;
      src12 <= 64'h74b7061c09ce15a8;
      src13 <= 64'h1eb95739b8acdd81;
      src14 <= 64'h7efa2faf58ba0bf3;
      src15 <= 64'h8c626a9fee4e6bc;
      src16 <= 64'h8429aeae877e5ea1;
      src17 <= 64'h402988fdf8cc3f3b;
      src18 <= 64'hecadbb86f16f1487;
      src19 <= 64'he642965cde386aeb;
      src20 <= 64'hf3ca5f6427fa8b8a;
      src21 <= 64'h52b049944b1dd9fd;
      src22 <= 64'hfccae6b86e566274;
      src23 <= 64'hc9d0a7f400425fc6;
      src24 <= 64'hb2975c6918ff358;
      src25 <= 64'h300a21879cb9f9aa;
      src26 <= 64'hefa2ce128c833848;
      src27 <= 64'h878f40ed2c805ac7;
      src28 <= 64'h94665d45284b7bcd;
      src29 <= 64'hc1378e75627b9de7;
      src30 <= 64'h4fb7c3bb4408c04c;
      src31 <= 64'hf23db30647caf779;
      src32 <= 64'hfd768f635163de1d;
      src33 <= 64'hcaa0a6796e83a7b2;
      src34 <= 64'h903374bfc81236e6;
      src35 <= 64'he65a3ae43a72017d;
      src36 <= 64'ha1832fdb31cb5e8e;
      src37 <= 64'hb3390a6ea0b87e45;
      src38 <= 64'h4643d7053df8eeef;
      src39 <= 64'hb47a5dcecf709452;
      src40 <= 64'h30331476f53fc3dd;
      src41 <= 64'hec6e61bd70c455a9;
      src42 <= 64'hf0bd7405650dd400;
      src43 <= 64'hc602bd20c1fa924e;
      src44 <= 64'h53e836639c14940d;
      src45 <= 64'h7b6e28f4e98ce25;
      src46 <= 64'hc334f55802cee581;
      src47 <= 64'hc329870a33e9e55e;
      src48 <= 64'h4741ee56b5e2834d;
      src49 <= 64'h6389bd3d26eeeba;
      src50 <= 64'haa5658322a5a421;
      src51 <= 64'hdd6d47e490e0172f;
      src52 <= 64'h12677895c6be596;
      src53 <= 64'hb7a02afd30d6863f;
      src54 <= 64'h8a663359abe0a177;
      src55 <= 64'h67fece7f1ff06dc;
      src56 <= 64'he7bf9a9664849eb5;
      src57 <= 64'h466bd06fa2b4d215;
      src58 <= 64'h82f1240d4e5c6dd2;
      src59 <= 64'he91e70af224af354;
      src60 <= 64'hb93c2989c399fd7f;
      src61 <= 64'hd020baee95fc7389;
      src62 <= 64'h8f4ed44214aaaefe;
      src63 <= 64'h43fd46ffd03459a4;
      #1
      src00 <= 64'h42ce91c0ccd9f2af;
      src01 <= 64'hb56b9357b34dc8b0;
      src02 <= 64'h1257363cf25dcb50;
      src03 <= 64'hca8033a7a5fd89c8;
      src04 <= 64'h85b303d3756b6c0d;
      src05 <= 64'h2287401ba7bbaa76;
      src06 <= 64'h8e50c79ac5826444;
      src07 <= 64'h57e7ef7b848610cf;
      src08 <= 64'hc65d8e4ed01e488b;
      src09 <= 64'h91fd7d4a5a31a6a6;
      src10 <= 64'hd560e64c55f7792a;
      src11 <= 64'h22d801701e6cbd83;
      src12 <= 64'h5d156b6eceec38d;
      src13 <= 64'h20068c1cbbd743b3;
      src14 <= 64'hb4cba0a317eeb1d;
      src15 <= 64'hcbf8e26a4fae667b;
      src16 <= 64'hed469bf4d5cf2dc4;
      src17 <= 64'hdd35d11688181a8;
      src18 <= 64'hc1a7de009ec12fa2;
      src19 <= 64'hcdc39412d95e17e1;
      src20 <= 64'h2e4025346987b052;
      src21 <= 64'hcd6a5e0c74279656;
      src22 <= 64'hf30459cc30c42d61;
      src23 <= 64'h5b8c4949106861d3;
      src24 <= 64'h6b42b6f1f94e3c8;
      src25 <= 64'h2d5590c905765983;
      src26 <= 64'h37e5725e5a1bdae;
      src27 <= 64'h79fe0a1b7efbe877;
      src28 <= 64'h1480f037d39a4bb0;
      src29 <= 64'hf484878d5bc9e889;
      src30 <= 64'hf7d870b678ac8704;
      src31 <= 64'hce03a34da022dfee;
      src32 <= 64'h96bfafff5b7751f;
      src33 <= 64'h5672ebc7606e8502;
      src34 <= 64'h291a58af259a2b28;
      src35 <= 64'hebbe1a41c781e11f;
      src36 <= 64'hae09ccfba3dee81f;
      src37 <= 64'hb4ea16d65ea29d1;
      src38 <= 64'ha2bb62833d83ad7c;
      src39 <= 64'h5a220eb23cf9d1fe;
      src40 <= 64'he0db22d329e316ad;
      src41 <= 64'h2353d45590bccb66;
      src42 <= 64'hc5507d2b909e7f78;
      src43 <= 64'hafdb4e0b01716f1d;
      src44 <= 64'hcd34bcd7b7ed75b4;
      src45 <= 64'h261cec19fff83cec;
      src46 <= 64'hd2f7442906714938;
      src47 <= 64'hf2460382951fe0;
      src48 <= 64'hc740525525cf51c4;
      src49 <= 64'hc96ef1a5ac707464;
      src50 <= 64'h6c4e109c9a6e611;
      src51 <= 64'hec2b5e213f7a38e0;
      src52 <= 64'h829fe7ba5d30db82;
      src53 <= 64'h667fceeb8889832c;
      src54 <= 64'h3ee29e686fa00319;
      src55 <= 64'hff7acd86409b3c5b;
      src56 <= 64'h86ce563de291f5e1;
      src57 <= 64'hc79385209c921e7f;
      src58 <= 64'h3cad275ae072caae;
      src59 <= 64'h9c684df10a515e87;
      src60 <= 64'hcc4e66dade0989b9;
      src61 <= 64'ha0483bb2f6d080c4;
      src62 <= 64'h64a2bc48f9fb4010;
      src63 <= 64'h9aabd22d75ef8aab;
      #1
      src00 <= 64'h2b6b7b4229502326;
      src01 <= 64'h693d993c796f9881;
      src02 <= 64'h586d7f415e47c2a0;
      src03 <= 64'hdccbbedc0e0d55b;
      src04 <= 64'hf5141524e08c28eb;
      src05 <= 64'h4bc972ce531da6ac;
      src06 <= 64'ha9d499ca2698c2d;
      src07 <= 64'h6e63ffa48d2ad974;
      src08 <= 64'h69199a8aaea62315;
      src09 <= 64'hba5612f7600aa45e;
      src10 <= 64'h22587c8958ccf9b4;
      src11 <= 64'h9cf600ec1c3c8d35;
      src12 <= 64'h7fe6a4e2a6f1e47;
      src13 <= 64'h65fd5f6993a25c9b;
      src14 <= 64'hae4a741ab5004950;
      src15 <= 64'h8dcd7d64b9e8e4ee;
      src16 <= 64'h2728ec952b52dab1;
      src17 <= 64'h3a6e8f122a1ace85;
      src18 <= 64'haf273f4055cdd72e;
      src19 <= 64'hd68d2bc2dac7c336;
      src20 <= 64'hdcfbde0ac5fee487;
      src21 <= 64'h2887a3a9e63317c3;
      src22 <= 64'he983cc1d25033a3e;
      src23 <= 64'h4e245cf78e33dcab;
      src24 <= 64'h58b5f05260e9bd79;
      src25 <= 64'hf6f259264e60678b;
      src26 <= 64'h25cc2478276d7e19;
      src27 <= 64'h8461f840e1a9344e;
      src28 <= 64'h1c769e1f83719849;
      src29 <= 64'h603803f32b2bcfda;
      src30 <= 64'h938ad77cb18d6a4;
      src31 <= 64'he47516941d8ac1a9;
      src32 <= 64'hb8f35c26d13ec39c;
      src33 <= 64'hec3826bc3a8d1c00;
      src34 <= 64'h2b02237ee2cd159a;
      src35 <= 64'h3544f189a9204633;
      src36 <= 64'haf04ef81b5481bf2;
      src37 <= 64'heb6ec9e0225f5457;
      src38 <= 64'he29b24d72bdc9c10;
      src39 <= 64'h55a3a12967ba6b1a;
      src40 <= 64'hdf98377981bd5336;
      src41 <= 64'h64e322cfa51de78b;
      src42 <= 64'h2e57386443eb280e;
      src43 <= 64'h5d4438218a7f03ae;
      src44 <= 64'heab3c4d8d4e4004b;
      src45 <= 64'h7a658abe1188afa1;
      src46 <= 64'hf3fa861390ed41f4;
      src47 <= 64'h179d221d8e5f37fa;
      src48 <= 64'h4bf41e101c622f82;
      src49 <= 64'hcfd645605c05c1f3;
      src50 <= 64'h1ce5fc632d116fe;
      src51 <= 64'hee65afeb1b674518;
      src52 <= 64'haf8c96a918f7e499;
      src53 <= 64'h3a05c0b73ddf55b2;
      src54 <= 64'hfbf70946d6ada066;
      src55 <= 64'h398071b14642cddb;
      src56 <= 64'h17776c3a57435d9c;
      src57 <= 64'h92dbd6134e051eea;
      src58 <= 64'hbd2cdb8d39ebfa32;
      src59 <= 64'h253df737c2185e77;
      src60 <= 64'hef96a21449b3fe66;
      src61 <= 64'hc6b7e7cbbe0d24ed;
      src62 <= 64'h486c0adf5bf26ec8;
      src63 <= 64'h1e94eb4bc74f73ca;
      #1
      src00 <= 64'h5bd71dc6ea75e34d;
      src01 <= 64'hfe38f4ebb6e0eac2;
      src02 <= 64'h1af4321addd3e779;
      src03 <= 64'h4a9686a4e7524102;
      src04 <= 64'h277dfc7b722c353d;
      src05 <= 64'h7fd2770a568d6f3e;
      src06 <= 64'hae5ceb3d1c275035;
      src07 <= 64'h6382f3b5f9adf8c5;
      src08 <= 64'hacf606fc387cdf02;
      src09 <= 64'h4fab2ad88091a21d;
      src10 <= 64'h6b8fd6af157ed9;
      src11 <= 64'h51306e5c78c5a976;
      src12 <= 64'hf325f875e4172ba3;
      src13 <= 64'hf7b37a86d21dbc09;
      src14 <= 64'ha5a0322c57842a9;
      src15 <= 64'h437249fd17ee2fe6;
      src16 <= 64'h53a9ec5db9b5c70e;
      src17 <= 64'h5d393bf9b2daa1f6;
      src18 <= 64'hf3f053233bd5f8a2;
      src19 <= 64'h213124bd01275a63;
      src20 <= 64'he998952cef58951f;
      src21 <= 64'hbdb62ff314e16706;
      src22 <= 64'hd9073286329cd43a;
      src23 <= 64'h6a4ace0ed89a9500;
      src24 <= 64'h61c61ae46a594b07;
      src25 <= 64'h183cfeceb09220;
      src26 <= 64'h44f20133f45c8840;
      src27 <= 64'hd3bb63d75e12425c;
      src28 <= 64'hb6ffe12c1a6f0c9a;
      src29 <= 64'h22ca9fe8a8aa7d13;
      src30 <= 64'h51cd2c07a8f78b61;
      src31 <= 64'h8f41d3e41eceb5e5;
      src32 <= 64'he93b4418b170b1ed;
      src33 <= 64'h7844c2ac729bd820;
      src34 <= 64'h8c3af69e74747f6f;
      src35 <= 64'h6a8d3e8420fe652b;
      src36 <= 64'hdcff697dd26d028d;
      src37 <= 64'h3f9bbcfc742c5905;
      src38 <= 64'h61f567969083bd6;
      src39 <= 64'he355c369b931a26d;
      src40 <= 64'hc67781b2c3a31607;
      src41 <= 64'h6df2fc823956fba9;
      src42 <= 64'h7a2be04940d2d16f;
      src43 <= 64'h3a6f36fa241813ef;
      src44 <= 64'h3006ff85166a1a98;
      src45 <= 64'h27b51ee70f1a6c44;
      src46 <= 64'hce1f40819f2d5db8;
      src47 <= 64'he668bb6ec408143f;
      src48 <= 64'had83095163eaa005;
      src49 <= 64'h7f00625769560c06;
      src50 <= 64'h64119d382ae201c0;
      src51 <= 64'hf60ce881c5ac7520;
      src52 <= 64'h855a7d8dd46e34aa;
      src53 <= 64'h53fb2ed1b9534807;
      src54 <= 64'h6f1d5baf952b750d;
      src55 <= 64'hedc641cd921bc646;
      src56 <= 64'h70fe3cfc991ab513;
      src57 <= 64'hd7f14ec29a9dadd2;
      src58 <= 64'hbb2966398e4a295d;
      src59 <= 64'hb2591c40021b632;
      src60 <= 64'h3e2b66532258edf3;
      src61 <= 64'h840658d1c1da8d39;
      src62 <= 64'h5690f74daedab7b5;
      src63 <= 64'h31307e46af797546;
      #1
      src00 <= 64'hb7ae77585b45cf5a;
      src01 <= 64'h77f4531bfde9d47d;
      src02 <= 64'hc06bad381d010478;
      src03 <= 64'hefb80c63f42f338f;
      src04 <= 64'hb44788bd5e2d2454;
      src05 <= 64'h67f8ab5705727bb5;
      src06 <= 64'hda98da57166adfc4;
      src07 <= 64'ha225183835e1392e;
      src08 <= 64'h7d5d9031e80bb7eb;
      src09 <= 64'hbb00d206f8542953;
      src10 <= 64'h3ea038fc095e099;
      src11 <= 64'h4fe4b7355c29b6da;
      src12 <= 64'hdd9539fcf7cd0b75;
      src13 <= 64'h5e15428a833cf90f;
      src14 <= 64'h42260a44773b8350;
      src15 <= 64'h72789d7597f0bfcf;
      src16 <= 64'h61f9c40838330558;
      src17 <= 64'hb44361f16c7354a;
      src18 <= 64'h7c2b940d9045a445;
      src19 <= 64'h6f48744f7abc9f0b;
      src20 <= 64'h1dd95d4c0637fdca;
      src21 <= 64'he299cb482449213a;
      src22 <= 64'hb49b93d51e709e19;
      src23 <= 64'h43a061c445a16970;
      src24 <= 64'h5804a8811d8cca3b;
      src25 <= 64'h39279358d5f52c0;
      src26 <= 64'h54e27ea64202faf9;
      src27 <= 64'h1152797ec20166e3;
      src28 <= 64'h20d5c16e961139cf;
      src29 <= 64'h393031a6c82a6c15;
      src30 <= 64'h3aeb5bc0f63d307c;
      src31 <= 64'h706146ffbecba4c8;
      src32 <= 64'he5039055f90b9724;
      src33 <= 64'h33672754da2e6e6c;
      src34 <= 64'hd4062cce773a13fb;
      src35 <= 64'h20e30a4dfbcefcd0;
      src36 <= 64'h1debf6c503ccb5;
      src37 <= 64'hd1bfbabaa908923b;
      src38 <= 64'hf33c4233c833b07e;
      src39 <= 64'hfaa2cbad467a6bdf;
      src40 <= 64'h8dff06d28340fed5;
      src41 <= 64'h72f78920dd7516f5;
      src42 <= 64'h68bfbf7ed4dc2301;
      src43 <= 64'hff28355076847398;
      src44 <= 64'h4bebcf4f2c94151d;
      src45 <= 64'h496749fbb2e02961;
      src46 <= 64'hd5e32aef05dd1ef0;
      src47 <= 64'hd87d3afca3705e8a;
      src48 <= 64'h5028361fa94501d7;
      src49 <= 64'h49954cf1faaf500c;
      src50 <= 64'hb55dc442c884e666;
      src51 <= 64'h23d83f2284403b37;
      src52 <= 64'h6b291a13637c3644;
      src53 <= 64'h39b66d71951a0518;
      src54 <= 64'h88653e42cefe73ec;
      src55 <= 64'h6c749cf41f7550bc;
      src56 <= 64'h854df9b62b66b1c0;
      src57 <= 64'h623a35ae7a31a27c;
      src58 <= 64'h14c30b503d0daad0;
      src59 <= 64'hd3100ac51932263c;
      src60 <= 64'h7ff5101d3f1cd31b;
      src61 <= 64'h677abeb744bfc434;
      src62 <= 64'hef05b6fed4879e7;
      src63 <= 64'h5b7801ea86343347;
   end
endmodule

