module compressor(
      input wire [127:0] src000,
      input wire [127:0] src001,
      input wire [127:0] src002,
      input wire [127:0] src003,
      input wire [127:0] src004,
      input wire [127:0] src005,
      input wire [127:0] src006,
      input wire [127:0] src007,
      input wire [127:0] src008,
      input wire [127:0] src009,
      input wire [127:0] src010,
      input wire [127:0] src011,
      input wire [127:0] src012,
      input wire [127:0] src013,
      input wire [127:0] src014,
      input wire [127:0] src015,
      input wire [127:0] src016,
      input wire [127:0] src017,
      input wire [127:0] src018,
      input wire [127:0] src019,
      input wire [127:0] src020,
      input wire [127:0] src021,
      input wire [127:0] src022,
      input wire [127:0] src023,
      input wire [127:0] src024,
      input wire [127:0] src025,
      input wire [127:0] src026,
      input wire [127:0] src027,
      input wire [127:0] src028,
      input wire [127:0] src029,
      input wire [127:0] src030,
      input wire [127:0] src031,
      input wire [127:0] src032,
      input wire [127:0] src033,
      input wire [127:0] src034,
      input wire [127:0] src035,
      input wire [127:0] src036,
      input wire [127:0] src037,
      input wire [127:0] src038,
      input wire [127:0] src039,
      input wire [127:0] src040,
      input wire [127:0] src041,
      input wire [127:0] src042,
      input wire [127:0] src043,
      input wire [127:0] src044,
      input wire [127:0] src045,
      input wire [127:0] src046,
      input wire [127:0] src047,
      input wire [127:0] src048,
      input wire [127:0] src049,
      input wire [127:0] src050,
      input wire [127:0] src051,
      input wire [127:0] src052,
      input wire [127:0] src053,
      input wire [127:0] src054,
      input wire [127:0] src055,
      input wire [127:0] src056,
      input wire [127:0] src057,
      input wire [127:0] src058,
      input wire [127:0] src059,
      input wire [127:0] src060,
      input wire [127:0] src061,
      input wire [127:0] src062,
      input wire [127:0] src063,
      input wire [127:0] src064,
      input wire [127:0] src065,
      input wire [127:0] src066,
      input wire [127:0] src067,
      input wire [127:0] src068,
      input wire [127:0] src069,
      input wire [127:0] src070,
      input wire [127:0] src071,
      input wire [127:0] src072,
      input wire [127:0] src073,
      input wire [127:0] src074,
      input wire [127:0] src075,
      input wire [127:0] src076,
      input wire [127:0] src077,
      input wire [127:0] src078,
      input wire [127:0] src079,
      input wire [127:0] src080,
      input wire [127:0] src081,
      input wire [127:0] src082,
      input wire [127:0] src083,
      input wire [127:0] src084,
      input wire [127:0] src085,
      input wire [127:0] src086,
      input wire [127:0] src087,
      input wire [127:0] src088,
      input wire [127:0] src089,
      input wire [127:0] src090,
      input wire [127:0] src091,
      input wire [127:0] src092,
      input wire [127:0] src093,
      input wire [127:0] src094,
      input wire [127:0] src095,
      input wire [127:0] src096,
      input wire [127:0] src097,
      input wire [127:0] src098,
      input wire [127:0] src099,
      input wire [127:0] src100,
      input wire [127:0] src101,
      input wire [127:0] src102,
      input wire [127:0] src103,
      input wire [127:0] src104,
      input wire [127:0] src105,
      input wire [127:0] src106,
      input wire [127:0] src107,
      input wire [127:0] src108,
      input wire [127:0] src109,
      input wire [127:0] src110,
      input wire [127:0] src111,
      input wire [127:0] src112,
      input wire [127:0] src113,
      input wire [127:0] src114,
      input wire [127:0] src115,
      input wire [127:0] src116,
      input wire [127:0] src117,
      input wire [127:0] src118,
      input wire [127:0] src119,
      input wire [127:0] src120,
      input wire [127:0] src121,
      input wire [127:0] src122,
      input wire [127:0] src123,
      input wire [127:0] src124,
      input wire [127:0] src125,
      input wire [127:0] src126,
      input wire [127:0] src127,
      output wire [1:0] dst000,
      output wire [1:0] dst001,
      output wire [1:0] dst002,
      output wire [0:0] dst003,
      output wire [0:0] dst004,
      output wire [1:0] dst005,
      output wire [0:0] dst006,
      output wire [1:0] dst007,
      output wire [1:0] dst008,
      output wire [1:0] dst009,
      output wire [1:0] dst010,
      output wire [1:0] dst011,
      output wire [1:0] dst012,
      output wire [0:0] dst013,
      output wire [1:0] dst014,
      output wire [1:0] dst015,
      output wire [1:0] dst016,
      output wire [1:0] dst017,
      output wire [1:0] dst018,
      output wire [1:0] dst019,
      output wire [1:0] dst020,
      output wire [1:0] dst021,
      output wire [1:0] dst022,
      output wire [1:0] dst023,
      output wire [1:0] dst024,
      output wire [1:0] dst025,
      output wire [1:0] dst026,
      output wire [1:0] dst027,
      output wire [1:0] dst028,
      output wire [1:0] dst029,
      output wire [1:0] dst030,
      output wire [1:0] dst031,
      output wire [1:0] dst032,
      output wire [1:0] dst033,
      output wire [1:0] dst034,
      output wire [1:0] dst035,
      output wire [1:0] dst036,
      output wire [1:0] dst037,
      output wire [0:0] dst038,
      output wire [0:0] dst039,
      output wire [1:0] dst040,
      output wire [1:0] dst041,
      output wire [1:0] dst042,
      output wire [1:0] dst043,
      output wire [1:0] dst044,
      output wire [1:0] dst045,
      output wire [1:0] dst046,
      output wire [1:0] dst047,
      output wire [1:0] dst048,
      output wire [1:0] dst049,
      output wire [1:0] dst050,
      output wire [1:0] dst051,
      output wire [1:0] dst052,
      output wire [1:0] dst053,
      output wire [1:0] dst054,
      output wire [1:0] dst055,
      output wire [1:0] dst056,
      output wire [1:0] dst057,
      output wire [1:0] dst058,
      output wire [1:0] dst059,
      output wire [1:0] dst060,
      output wire [0:0] dst061,
      output wire [1:0] dst062,
      output wire [1:0] dst063,
      output wire [1:0] dst064,
      output wire [1:0] dst065,
      output wire [1:0] dst066,
      output wire [0:0] dst067,
      output wire [1:0] dst068,
      output wire [1:0] dst069,
      output wire [1:0] dst070,
      output wire [1:0] dst071,
      output wire [1:0] dst072,
      output wire [1:0] dst073,
      output wire [1:0] dst074,
      output wire [1:0] dst075,
      output wire [1:0] dst076,
      output wire [1:0] dst077,
      output wire [1:0] dst078,
      output wire [1:0] dst079,
      output wire [1:0] dst080,
      output wire [1:0] dst081,
      output wire [1:0] dst082,
      output wire [0:0] dst083,
      output wire [1:0] dst084,
      output wire [1:0] dst085,
      output wire [1:0] dst086,
      output wire [1:0] dst087,
      output wire [1:0] dst088,
      output wire [1:0] dst089,
      output wire [1:0] dst090,
      output wire [1:0] dst091,
      output wire [1:0] dst092,
      output wire [1:0] dst093,
      output wire [1:0] dst094,
      output wire [1:0] dst095,
      output wire [1:0] dst096,
      output wire [1:0] dst097,
      output wire [1:0] dst098,
      output wire [1:0] dst099,
      output wire [1:0] dst100,
      output wire [1:0] dst101,
      output wire [1:0] dst102,
      output wire [1:0] dst103,
      output wire [1:0] dst104,
      output wire [1:0] dst105,
      output wire [1:0] dst106,
      output wire [1:0] dst107,
      output wire [1:0] dst108,
      output wire [1:0] dst109,
      output wire [1:0] dst110,
      output wire [1:0] dst111,
      output wire [0:0] dst112,
      output wire [1:0] dst113,
      output wire [1:0] dst114,
      output wire [1:0] dst115,
      output wire [1:0] dst116,
      output wire [1:0] dst117,
      output wire [1:0] dst118,
      output wire [1:0] dst119,
      output wire [1:0] dst120,
      output wire [0:0] dst121,
      output wire [1:0] dst122,
      output wire [1:0] dst123,
      output wire [1:0] dst124,
      output wire [1:0] dst125,
      output wire [1:0] dst126,
      output wire [1:0] dst127,
      output wire [1:0] dst128,
      output wire [1:0] dst129,
      output wire [1:0] dst130,
      output wire [1:0] dst131,
      output wire [1:0] dst132,
      output wire [1:0] dst133,
      output wire [0:0] dst134
   );
   wire [193:0] stage000;
   wire [231:0] stage001;
   wire [247:0] stage002;
   wire [219:0] stage003;
   wire [277:0] stage004;
   wire [283:0] stage005;
   wire [260:0] stage006;
   wire [261:0] stage007;
   wire [249:0] stage008;
   wire [245:0] stage009;
   wire [302:0] stage010;
   wire [267:0] stage011;
   wire [328:0] stage012;
   wire [274:0] stage013;
   wire [310:0] stage014;
   wire [264:0] stage015;
   wire [294:0] stage016;
   wire [287:0] stage017;
   wire [257:0] stage018;
   wire [281:0] stage019;
   wire [237:0] stage020;
   wire [302:0] stage021;
   wire [236:0] stage022;
   wire [321:0] stage023;
   wire [262:0] stage024;
   wire [303:0] stage025;
   wire [248:0] stage026;
   wire [242:0] stage027;
   wire [273:0] stage028;
   wire [294:0] stage029;
   wire [250:0] stage030;
   wire [258:0] stage031;
   wire [308:0] stage032;
   wire [304:0] stage033;
   wire [315:0] stage034;
   wire [269:0] stage035;
   wire [234:0] stage036;
   wire [283:0] stage037;
   wire [261:0] stage038;
   wire [259:0] stage039;
   wire [310:0] stage040;
   wire [286:0] stage041;
   wire [300:0] stage042;
   wire [224:0] stage043;
   wire [232:0] stage044;
   wire [277:0] stage045;
   wire [282:0] stage046;
   wire [240:0] stage047;
   wire [350:0] stage048;
   wire [262:0] stage049;
   wire [288:0] stage050;
   wire [262:0] stage051;
   wire [283:0] stage052;
   wire [257:0] stage053;
   wire [265:0] stage054;
   wire [303:0] stage055;
   wire [296:0] stage056;
   wire [263:0] stage057;
   wire [240:0] stage058;
   wire [325:0] stage059;
   wire [253:0] stage060;
   wire [283:0] stage061;
   wire [262:0] stage062;
   wire [226:0] stage063;
   wire [272:0] stage064;
   wire [269:0] stage065;
   wire [292:0] stage066;
   wire [270:0] stage067;
   wire [288:0] stage068;
   wire [277:0] stage069;
   wire [269:0] stage070;
   wire [271:0] stage071;
   wire [317:0] stage072;
   wire [252:0] stage073;
   wire [267:0] stage074;
   wire [215:0] stage075;
   wire [221:0] stage076;
   wire [270:0] stage077;
   wire [239:0] stage078;
   wire [264:0] stage079;
   wire [269:0] stage080;
   wire [299:0] stage081;
   wire [272:0] stage082;
   wire [282:0] stage083;
   wire [249:0] stage084;
   wire [280:0] stage085;
   wire [297:0] stage086;
   wire [245:0] stage087;
   wire [287:0] stage088;
   wire [277:0] stage089;
   wire [260:0] stage090;
   wire [345:0] stage091;
   wire [259:0] stage092;
   wire [242:0] stage093;
   wire [251:0] stage094;
   wire [231:0] stage095;
   wire [248:0] stage096;
   wire [234:0] stage097;
   wire [246:0] stage098;
   wire [304:0] stage099;
   wire [231:0] stage100;
   wire [272:0] stage101;
   wire [252:0] stage102;
   wire [262:0] stage103;
   wire [267:0] stage104;
   wire [231:0] stage105;
   wire [261:0] stage106;
   wire [268:0] stage107;
   wire [265:0] stage108;
   wire [237:0] stage109;
   wire [273:0] stage110;
   wire [266:0] stage111;
   wire [244:0] stage112;
   wire [243:0] stage113;
   wire [254:0] stage114;
   wire [264:0] stage115;
   wire [244:0] stage116;
   wire [265:0] stage117;
   wire [265:0] stage118;
   wire [242:0] stage119;
   wire [257:0] stage120;
   wire [241:0] stage121;
   wire [250:0] stage122;
   wire [329:0] stage123;
   wire [240:0] stage124;
   wire [287:0] stage125;
   wire [288:0] stage126;
   wire [292:0] stage127;
   wire [91:0] stage128;
   wire [87:0] stage129;
   wire [21:0] stage130;
   wire [17:0] stage131;
   wire [8:0] stage132;
   wire [7:0] stage133;
   wire [0:0] stage134;
   assign stage000[127:0] = src000;
   assign stage001[127:0] = src001;
   assign stage002[127:0] = src002;
   assign stage003[127:0] = src003;
   assign stage004[127:0] = src004;
   assign stage005[127:0] = src005;
   assign stage006[127:0] = src006;
   assign stage007[127:0] = src007;
   assign stage008[127:0] = src008;
   assign stage009[127:0] = src009;
   assign stage010[127:0] = src010;
   assign stage011[127:0] = src011;
   assign stage012[127:0] = src012;
   assign stage013[127:0] = src013;
   assign stage014[127:0] = src014;
   assign stage015[127:0] = src015;
   assign stage016[127:0] = src016;
   assign stage017[127:0] = src017;
   assign stage018[127:0] = src018;
   assign stage019[127:0] = src019;
   assign stage020[127:0] = src020;
   assign stage021[127:0] = src021;
   assign stage022[127:0] = src022;
   assign stage023[127:0] = src023;
   assign stage024[127:0] = src024;
   assign stage025[127:0] = src025;
   assign stage026[127:0] = src026;
   assign stage027[127:0] = src027;
   assign stage028[127:0] = src028;
   assign stage029[127:0] = src029;
   assign stage030[127:0] = src030;
   assign stage031[127:0] = src031;
   assign stage032[127:0] = src032;
   assign stage033[127:0] = src033;
   assign stage034[127:0] = src034;
   assign stage035[127:0] = src035;
   assign stage036[127:0] = src036;
   assign stage037[127:0] = src037;
   assign stage038[127:0] = src038;
   assign stage039[127:0] = src039;
   assign stage040[127:0] = src040;
   assign stage041[127:0] = src041;
   assign stage042[127:0] = src042;
   assign stage043[127:0] = src043;
   assign stage044[127:0] = src044;
   assign stage045[127:0] = src045;
   assign stage046[127:0] = src046;
   assign stage047[127:0] = src047;
   assign stage048[127:0] = src048;
   assign stage049[127:0] = src049;
   assign stage050[127:0] = src050;
   assign stage051[127:0] = src051;
   assign stage052[127:0] = src052;
   assign stage053[127:0] = src053;
   assign stage054[127:0] = src054;
   assign stage055[127:0] = src055;
   assign stage056[127:0] = src056;
   assign stage057[127:0] = src057;
   assign stage058[127:0] = src058;
   assign stage059[127:0] = src059;
   assign stage060[127:0] = src060;
   assign stage061[127:0] = src061;
   assign stage062[127:0] = src062;
   assign stage063[127:0] = src063;
   assign stage064[127:0] = src064;
   assign stage065[127:0] = src065;
   assign stage066[127:0] = src066;
   assign stage067[127:0] = src067;
   assign stage068[127:0] = src068;
   assign stage069[127:0] = src069;
   assign stage070[127:0] = src070;
   assign stage071[127:0] = src071;
   assign stage072[127:0] = src072;
   assign stage073[127:0] = src073;
   assign stage074[127:0] = src074;
   assign stage075[127:0] = src075;
   assign stage076[127:0] = src076;
   assign stage077[127:0] = src077;
   assign stage078[127:0] = src078;
   assign stage079[127:0] = src079;
   assign stage080[127:0] = src080;
   assign stage081[127:0] = src081;
   assign stage082[127:0] = src082;
   assign stage083[127:0] = src083;
   assign stage084[127:0] = src084;
   assign stage085[127:0] = src085;
   assign stage086[127:0] = src086;
   assign stage087[127:0] = src087;
   assign stage088[127:0] = src088;
   assign stage089[127:0] = src089;
   assign stage090[127:0] = src090;
   assign stage091[127:0] = src091;
   assign stage092[127:0] = src092;
   assign stage093[127:0] = src093;
   assign stage094[127:0] = src094;
   assign stage095[127:0] = src095;
   assign stage096[127:0] = src096;
   assign stage097[127:0] = src097;
   assign stage098[127:0] = src098;
   assign stage099[127:0] = src099;
   assign stage100[127:0] = src100;
   assign stage101[127:0] = src101;
   assign stage102[127:0] = src102;
   assign stage103[127:0] = src103;
   assign stage104[127:0] = src104;
   assign stage105[127:0] = src105;
   assign stage106[127:0] = src106;
   assign stage107[127:0] = src107;
   assign stage108[127:0] = src108;
   assign stage109[127:0] = src109;
   assign stage110[127:0] = src110;
   assign stage111[127:0] = src111;
   assign stage112[127:0] = src112;
   assign stage113[127:0] = src113;
   assign stage114[127:0] = src114;
   assign stage115[127:0] = src115;
   assign stage116[127:0] = src116;
   assign stage117[127:0] = src117;
   assign stage118[127:0] = src118;
   assign stage119[127:0] = src119;
   assign stage120[127:0] = src120;
   assign stage121[127:0] = src121;
   assign stage122[127:0] = src122;
   assign stage123[127:0] = src123;
   assign stage124[127:0] = src124;
   assign stage125[127:0] = src125;
   assign stage126[127:0] = src126;
   assign stage127[127:0] = src127;
   assign dst000 = stage000[193:192];
   assign dst001 = stage001[231:230];
   assign dst002 = stage002[247:246];
   assign dst003 = stage003[219:219];
   assign dst004 = stage004[277:277];
   assign dst005 = stage005[283:282];
   assign dst006 = stage006[260:260];
   assign dst007 = stage007[261:260];
   assign dst008 = stage008[249:248];
   assign dst009 = stage009[245:244];
   assign dst010 = stage010[302:301];
   assign dst011 = stage011[267:266];
   assign dst012 = stage012[328:327];
   assign dst013 = stage013[274:274];
   assign dst014 = stage014[310:309];
   assign dst015 = stage015[264:263];
   assign dst016 = stage016[294:293];
   assign dst017 = stage017[287:286];
   assign dst018 = stage018[257:256];
   assign dst019 = stage019[281:280];
   assign dst020 = stage020[237:236];
   assign dst021 = stage021[302:301];
   assign dst022 = stage022[236:235];
   assign dst023 = stage023[321:320];
   assign dst024 = stage024[262:261];
   assign dst025 = stage025[303:302];
   assign dst026 = stage026[248:247];
   assign dst027 = stage027[242:241];
   assign dst028 = stage028[273:272];
   assign dst029 = stage029[294:293];
   assign dst030 = stage030[250:249];
   assign dst031 = stage031[258:257];
   assign dst032 = stage032[308:307];
   assign dst033 = stage033[304:303];
   assign dst034 = stage034[315:314];
   assign dst035 = stage035[269:268];
   assign dst036 = stage036[234:233];
   assign dst037 = stage037[283:282];
   assign dst038 = stage038[261:261];
   assign dst039 = stage039[259:259];
   assign dst040 = stage040[310:309];
   assign dst041 = stage041[286:285];
   assign dst042 = stage042[300:299];
   assign dst043 = stage043[224:223];
   assign dst044 = stage044[232:231];
   assign dst045 = stage045[277:276];
   assign dst046 = stage046[282:281];
   assign dst047 = stage047[240:239];
   assign dst048 = stage048[350:349];
   assign dst049 = stage049[262:261];
   assign dst050 = stage050[288:287];
   assign dst051 = stage051[262:261];
   assign dst052 = stage052[283:282];
   assign dst053 = stage053[257:256];
   assign dst054 = stage054[265:264];
   assign dst055 = stage055[303:302];
   assign dst056 = stage056[296:295];
   assign dst057 = stage057[263:262];
   assign dst058 = stage058[240:239];
   assign dst059 = stage059[325:324];
   assign dst060 = stage060[253:252];
   assign dst061 = stage061[283:283];
   assign dst062 = stage062[262:261];
   assign dst063 = stage063[226:225];
   assign dst064 = stage064[272:271];
   assign dst065 = stage065[269:268];
   assign dst066 = stage066[292:291];
   assign dst067 = stage067[270:270];
   assign dst068 = stage068[288:287];
   assign dst069 = stage069[277:276];
   assign dst070 = stage070[269:268];
   assign dst071 = stage071[271:270];
   assign dst072 = stage072[317:316];
   assign dst073 = stage073[252:251];
   assign dst074 = stage074[267:266];
   assign dst075 = stage075[215:214];
   assign dst076 = stage076[221:220];
   assign dst077 = stage077[270:269];
   assign dst078 = stage078[239:238];
   assign dst079 = stage079[264:263];
   assign dst080 = stage080[269:268];
   assign dst081 = stage081[299:298];
   assign dst082 = stage082[272:271];
   assign dst083 = stage083[282:282];
   assign dst084 = stage084[249:248];
   assign dst085 = stage085[280:279];
   assign dst086 = stage086[297:296];
   assign dst087 = stage087[245:244];
   assign dst088 = stage088[287:286];
   assign dst089 = stage089[277:276];
   assign dst090 = stage090[260:259];
   assign dst091 = stage091[345:344];
   assign dst092 = stage092[259:258];
   assign dst093 = stage093[242:241];
   assign dst094 = stage094[251:250];
   assign dst095 = stage095[231:230];
   assign dst096 = stage096[248:247];
   assign dst097 = stage097[234:233];
   assign dst098 = stage098[246:245];
   assign dst099 = stage099[304:303];
   assign dst100 = stage100[231:230];
   assign dst101 = stage101[272:271];
   assign dst102 = stage102[252:251];
   assign dst103 = stage103[262:261];
   assign dst104 = stage104[267:266];
   assign dst105 = stage105[231:230];
   assign dst106 = stage106[261:260];
   assign dst107 = stage107[268:267];
   assign dst108 = stage108[265:264];
   assign dst109 = stage109[237:236];
   assign dst110 = stage110[273:272];
   assign dst111 = stage111[266:265];
   assign dst112 = stage112[244:244];
   assign dst113 = stage113[243:242];
   assign dst114 = stage114[254:253];
   assign dst115 = stage115[264:263];
   assign dst116 = stage116[244:243];
   assign dst117 = stage117[265:264];
   assign dst118 = stage118[265:264];
   assign dst119 = stage119[242:241];
   assign dst120 = stage120[257:256];
   assign dst121 = stage121[241:241];
   assign dst122 = stage122[250:249];
   assign dst123 = stage123[329:328];
   assign dst124 = stage124[240:239];
   assign dst125 = stage125[287:286];
   assign dst126 = stage126[288:287];
   assign dst127 = stage127[292:291];
   assign dst128 = stage128[91:90];
   assign dst129 = stage129[87:86];
   assign dst130 = stage130[21:20];
   assign dst131 = stage131[17:16];
   assign dst132 = stage132[8:7];
   assign dst133 = stage133[7:6];
   assign dst134 = stage134[0:0];
   gpc1_1 gpc1_1_0(
      {stage000[0]},
      {stage000[128]}
   );
   gpc1_1 gpc1_1_1(
      {stage000[1]},
      {stage000[129]}
   );
   gpc1_1 gpc1_1_2(
      {stage000[2]},
      {stage000[130]}
   );
   gpc1_1 gpc1_1_3(
      {stage000[3]},
      {stage000[131]}
   );
   gpc1_1 gpc1_1_4(
      {stage000[4]},
      {stage000[132]}
   );
   gpc1_1 gpc1_1_5(
      {stage000[5]},
      {stage000[133]}
   );
   gpc1_1 gpc1_1_6(
      {stage000[6]},
      {stage000[134]}
   );
   gpc1_1 gpc1_1_7(
      {stage000[7]},
      {stage000[135]}
   );
   gpc1_1 gpc1_1_8(
      {stage000[8]},
      {stage000[136]}
   );
   gpc1_1 gpc1_1_9(
      {stage000[9]},
      {stage000[137]}
   );
   gpc1_1 gpc1_1_10(
      {stage000[10]},
      {stage000[138]}
   );
   gpc1_1 gpc1_1_11(
      {stage000[11]},
      {stage000[139]}
   );
   gpc1_1 gpc1_1_12(
      {stage000[12]},
      {stage000[140]}
   );
   gpc1_1 gpc1_1_13(
      {stage000[13]},
      {stage000[141]}
   );
   gpc1_1 gpc1_1_14(
      {stage000[14]},
      {stage000[142]}
   );
   gpc1_1 gpc1_1_15(
      {stage000[15]},
      {stage000[143]}
   );
   gpc1_1 gpc1_1_16(
      {stage000[16]},
      {stage000[144]}
   );
   gpc1_1 gpc1_1_17(
      {stage000[17]},
      {stage000[145]}
   );
   gpc1_1 gpc1_1_18(
      {stage000[18]},
      {stage000[146]}
   );
   gpc1_1 gpc1_1_19(
      {stage000[19]},
      {stage000[147]}
   );
   gpc1_1 gpc1_1_20(
      {stage000[20]},
      {stage000[148]}
   );
   gpc606_5 gpc606_5_21(
      {stage000[21], stage000[22], stage000[23], stage000[24], stage000[25], stage000[26]},
      {stage002[0], stage002[1], stage002[2], stage002[3], stage002[4], stage002[5]},
      {stage004[128], stage003[128], stage002[128], stage001[128], stage000[149]}
   );
   gpc606_5 gpc606_5_22(
      {stage000[27], stage000[28], stage000[29], stage000[30], stage000[31], stage000[32]},
      {stage002[6], stage002[7], stage002[8], stage002[9], stage002[10], stage002[11]},
      {stage004[129], stage003[129], stage002[129], stage001[129], stage000[150]}
   );
   gpc615_5 gpc615_5_23(
      {stage000[33], stage000[34], stage000[35], stage000[36], stage000[37]},
      {stage001[0]},
      {stage002[12], stage002[13], stage002[14], stage002[15], stage002[16], stage002[17]},
      {stage004[130], stage003[130], stage002[130], stage001[130], stage000[151]}
   );
   gpc615_5 gpc615_5_24(
      {stage000[38], stage000[39], stage000[40], stage000[41], stage000[42]},
      {stage001[1]},
      {stage002[18], stage002[19], stage002[20], stage002[21], stage002[22], stage002[23]},
      {stage004[131], stage003[131], stage002[131], stage001[131], stage000[152]}
   );
   gpc615_5 gpc615_5_25(
      {stage000[43], stage000[44], stage000[45], stage000[46], stage000[47]},
      {stage001[2]},
      {stage002[24], stage002[25], stage002[26], stage002[27], stage002[28], stage002[29]},
      {stage004[132], stage003[132], stage002[132], stage001[132], stage000[153]}
   );
   gpc615_5 gpc615_5_26(
      {stage000[48], stage000[49], stage000[50], stage000[51], stage000[52]},
      {stage001[3]},
      {stage002[30], stage002[31], stage002[32], stage002[33], stage002[34], stage002[35]},
      {stage004[133], stage003[133], stage002[133], stage001[133], stage000[154]}
   );
   gpc2135_5 gpc2135_5_27(
      {stage000[53], stage000[54], stage000[55], stage000[56], stage000[57]},
      {stage001[4], stage001[5], stage001[6]},
      {stage002[36]},
      {stage003[0], stage003[1]},
      {stage004[134], stage003[134], stage002[134], stage001[134], stage000[155]}
   );
   gpc2135_5 gpc2135_5_28(
      {stage000[58], stage000[59], stage000[60], stage000[61], stage000[62]},
      {stage001[7], stage001[8], stage001[9]},
      {stage002[37]},
      {stage003[2], stage003[3]},
      {stage004[135], stage003[135], stage002[135], stage001[135], stage000[156]}
   );
   gpc2135_5 gpc2135_5_29(
      {stage000[63], stage000[64], stage000[65], stage000[66], stage000[67]},
      {stage001[10], stage001[11], stage001[12]},
      {stage002[38]},
      {stage003[4], stage003[5]},
      {stage004[136], stage003[136], stage002[136], stage001[136], stage000[157]}
   );
   gpc2135_5 gpc2135_5_30(
      {stage000[68], stage000[69], stage000[70], stage000[71], stage000[72]},
      {stage001[13], stage001[14], stage001[15]},
      {stage002[39]},
      {stage003[6], stage003[7]},
      {stage004[137], stage003[137], stage002[137], stage001[137], stage000[158]}
   );
   gpc2135_5 gpc2135_5_31(
      {stage000[73], stage000[74], stage000[75], stage000[76], stage000[77]},
      {stage001[16], stage001[17], stage001[18]},
      {stage002[40]},
      {stage003[8], stage003[9]},
      {stage004[138], stage003[138], stage002[138], stage001[138], stage000[159]}
   );
   gpc2135_5 gpc2135_5_32(
      {stage000[78], stage000[79], stage000[80], stage000[81], stage000[82]},
      {stage001[19], stage001[20], stage001[21]},
      {stage002[41]},
      {stage003[10], stage003[11]},
      {stage004[139], stage003[139], stage002[139], stage001[139], stage000[160]}
   );
   gpc2135_5 gpc2135_5_33(
      {stage000[83], stage000[84], stage000[85], stage000[86], stage000[87]},
      {stage001[22], stage001[23], stage001[24]},
      {stage002[42]},
      {stage003[12], stage003[13]},
      {stage004[140], stage003[140], stage002[140], stage001[140], stage000[161]}
   );
   gpc2135_5 gpc2135_5_34(
      {stage000[88], stage000[89], stage000[90], stage000[91], stage000[92]},
      {stage001[25], stage001[26], stage001[27]},
      {stage002[43]},
      {stage003[14], stage003[15]},
      {stage004[141], stage003[141], stage002[141], stage001[141], stage000[162]}
   );
   gpc2135_5 gpc2135_5_35(
      {stage000[93], stage000[94], stage000[95], stage000[96], stage000[97]},
      {stage001[28], stage001[29], stage001[30]},
      {stage002[44]},
      {stage003[16], stage003[17]},
      {stage004[142], stage003[142], stage002[142], stage001[142], stage000[163]}
   );
   gpc2135_5 gpc2135_5_36(
      {stage000[98], stage000[99], stage000[100], stage000[101], stage000[102]},
      {stage001[31], stage001[32], stage001[33]},
      {stage002[45]},
      {stage003[18], stage003[19]},
      {stage004[143], stage003[143], stage002[143], stage001[143], stage000[164]}
   );
   gpc2135_5 gpc2135_5_37(
      {stage000[103], stage000[104], stage000[105], stage000[106], stage000[107]},
      {stage001[34], stage001[35], stage001[36]},
      {stage002[46]},
      {stage003[20], stage003[21]},
      {stage004[144], stage003[144], stage002[144], stage001[144], stage000[165]}
   );
   gpc2135_5 gpc2135_5_38(
      {stage000[108], stage000[109], stage000[110], stage000[111], stage000[112]},
      {stage001[37], stage001[38], stage001[39]},
      {stage002[47]},
      {stage003[22], stage003[23]},
      {stage004[145], stage003[145], stage002[145], stage001[145], stage000[166]}
   );
   gpc2135_5 gpc2135_5_39(
      {stage000[113], stage000[114], stage000[115], stage000[116], stage000[117]},
      {stage001[40], stage001[41], stage001[42]},
      {stage002[48]},
      {stage003[24], stage003[25]},
      {stage004[146], stage003[146], stage002[146], stage001[146], stage000[167]}
   );
   gpc2135_5 gpc2135_5_40(
      {stage000[118], stage000[119], stage000[120], stage000[121], stage000[122]},
      {stage001[43], stage001[44], stage001[45]},
      {stage002[49]},
      {stage003[26], stage003[27]},
      {stage004[147], stage003[147], stage002[147], stage001[147], stage000[168]}
   );
   gpc2135_5 gpc2135_5_41(
      {stage000[123], stage000[124], stage000[125], stage000[126], stage000[127]},
      {stage001[46], stage001[47], stage001[48]},
      {stage002[50]},
      {stage003[28], stage003[29]},
      {stage004[148], stage003[148], stage002[148], stage001[148], stage000[169]}
   );
   gpc1_1 gpc1_1_42(
      {stage001[49]},
      {stage001[149]}
   );
   gpc1_1 gpc1_1_43(
      {stage001[50]},
      {stage001[150]}
   );
   gpc1_1 gpc1_1_44(
      {stage001[51]},
      {stage001[151]}
   );
   gpc1_1 gpc1_1_45(
      {stage001[52]},
      {stage001[152]}
   );
   gpc1_1 gpc1_1_46(
      {stage001[53]},
      {stage001[153]}
   );
   gpc1_1 gpc1_1_47(
      {stage001[54]},
      {stage001[154]}
   );
   gpc1_1 gpc1_1_48(
      {stage001[55]},
      {stage001[155]}
   );
   gpc1_1 gpc1_1_49(
      {stage001[56]},
      {stage001[156]}
   );
   gpc1_1 gpc1_1_50(
      {stage001[57]},
      {stage001[157]}
   );
   gpc1_1 gpc1_1_51(
      {stage001[58]},
      {stage001[158]}
   );
   gpc1_1 gpc1_1_52(
      {stage001[59]},
      {stage001[159]}
   );
   gpc1_1 gpc1_1_53(
      {stage001[60]},
      {stage001[160]}
   );
   gpc1_1 gpc1_1_54(
      {stage001[61]},
      {stage001[161]}
   );
   gpc1_1 gpc1_1_55(
      {stage001[62]},
      {stage001[162]}
   );
   gpc1_1 gpc1_1_56(
      {stage001[63]},
      {stage001[163]}
   );
   gpc1_1 gpc1_1_57(
      {stage001[64]},
      {stage001[164]}
   );
   gpc1_1 gpc1_1_58(
      {stage001[65]},
      {stage001[165]}
   );
   gpc1_1 gpc1_1_59(
      {stage001[66]},
      {stage001[166]}
   );
   gpc1_1 gpc1_1_60(
      {stage001[67]},
      {stage001[167]}
   );
   gpc1_1 gpc1_1_61(
      {stage001[68]},
      {stage001[168]}
   );
   gpc1_1 gpc1_1_62(
      {stage001[69]},
      {stage001[169]}
   );
   gpc1_1 gpc1_1_63(
      {stage001[70]},
      {stage001[170]}
   );
   gpc1_1 gpc1_1_64(
      {stage001[71]},
      {stage001[171]}
   );
   gpc1_1 gpc1_1_65(
      {stage001[72]},
      {stage001[172]}
   );
   gpc1_1 gpc1_1_66(
      {stage001[73]},
      {stage001[173]}
   );
   gpc606_5 gpc606_5_67(
      {stage001[74], stage001[75], stage001[76], stage001[77], stage001[78], stage001[79]},
      {stage003[30], stage003[31], stage003[32], stage003[33], stage003[34], stage003[35]},
      {stage005[128], stage004[149], stage003[149], stage002[149], stage001[174]}
   );
   gpc606_5 gpc606_5_68(
      {stage001[80], stage001[81], stage001[82], stage001[83], stage001[84], stage001[85]},
      {stage003[36], stage003[37], stage003[38], stage003[39], stage003[40], stage003[41]},
      {stage005[129], stage004[150], stage003[150], stage002[150], stage001[175]}
   );
   gpc606_5 gpc606_5_69(
      {stage001[86], stage001[87], stage001[88], stage001[89], stage001[90], stage001[91]},
      {stage003[42], stage003[43], stage003[44], stage003[45], stage003[46], stage003[47]},
      {stage005[130], stage004[151], stage003[151], stage002[151], stage001[176]}
   );
   gpc606_5 gpc606_5_70(
      {stage001[92], stage001[93], stage001[94], stage001[95], stage001[96], stage001[97]},
      {stage003[48], stage003[49], stage003[50], stage003[51], stage003[52], stage003[53]},
      {stage005[131], stage004[152], stage003[152], stage002[152], stage001[177]}
   );
   gpc606_5 gpc606_5_71(
      {stage001[98], stage001[99], stage001[100], stage001[101], stage001[102], stage001[103]},
      {stage003[54], stage003[55], stage003[56], stage003[57], stage003[58], stage003[59]},
      {stage005[132], stage004[153], stage003[153], stage002[153], stage001[178]}
   );
   gpc606_5 gpc606_5_72(
      {stage001[104], stage001[105], stage001[106], stage001[107], stage001[108], stage001[109]},
      {stage003[60], stage003[61], stage003[62], stage003[63], stage003[64], stage003[65]},
      {stage005[133], stage004[154], stage003[154], stage002[154], stage001[179]}
   );
   gpc606_5 gpc606_5_73(
      {stage001[110], stage001[111], stage001[112], stage001[113], stage001[114], stage001[115]},
      {stage003[66], stage003[67], stage003[68], stage003[69], stage003[70], stage003[71]},
      {stage005[134], stage004[155], stage003[155], stage002[155], stage001[180]}
   );
   gpc606_5 gpc606_5_74(
      {stage001[116], stage001[117], stage001[118], stage001[119], stage001[120], stage001[121]},
      {stage003[72], stage003[73], stage003[74], stage003[75], stage003[76], stage003[77]},
      {stage005[135], stage004[156], stage003[156], stage002[156], stage001[181]}
   );
   gpc606_5 gpc606_5_75(
      {stage001[122], stage001[123], stage001[124], stage001[125], stage001[126], stage001[127]},
      {stage003[78], stage003[79], stage003[80], stage003[81], stage003[82], stage003[83]},
      {stage005[136], stage004[157], stage003[157], stage002[157], stage001[182]}
   );
   gpc1_1 gpc1_1_76(
      {stage002[51]},
      {stage002[158]}
   );
   gpc1_1 gpc1_1_77(
      {stage002[52]},
      {stage002[159]}
   );
   gpc1_1 gpc1_1_78(
      {stage002[53]},
      {stage002[160]}
   );
   gpc1_1 gpc1_1_79(
      {stage002[54]},
      {stage002[161]}
   );
   gpc1_1 gpc1_1_80(
      {stage002[55]},
      {stage002[162]}
   );
   gpc1_1 gpc1_1_81(
      {stage002[56]},
      {stage002[163]}
   );
   gpc1_1 gpc1_1_82(
      {stage002[57]},
      {stage002[164]}
   );
   gpc1_1 gpc1_1_83(
      {stage002[58]},
      {stage002[165]}
   );
   gpc1_1 gpc1_1_84(
      {stage002[59]},
      {stage002[166]}
   );
   gpc1_1 gpc1_1_85(
      {stage002[60]},
      {stage002[167]}
   );
   gpc1_1 gpc1_1_86(
      {stage002[61]},
      {stage002[168]}
   );
   gpc1_1 gpc1_1_87(
      {stage002[62]},
      {stage002[169]}
   );
   gpc1_1 gpc1_1_88(
      {stage002[63]},
      {stage002[170]}
   );
   gpc1_1 gpc1_1_89(
      {stage002[64]},
      {stage002[171]}
   );
   gpc1_1 gpc1_1_90(
      {stage002[65]},
      {stage002[172]}
   );
   gpc1_1 gpc1_1_91(
      {stage002[66]},
      {stage002[173]}
   );
   gpc1_1 gpc1_1_92(
      {stage002[67]},
      {stage002[174]}
   );
   gpc1_1 gpc1_1_93(
      {stage002[68]},
      {stage002[175]}
   );
   gpc1_1 gpc1_1_94(
      {stage002[69]},
      {stage002[176]}
   );
   gpc1_1 gpc1_1_95(
      {stage002[70]},
      {stage002[177]}
   );
   gpc606_5 gpc606_5_96(
      {stage002[71], stage002[72], stage002[73], stage002[74], stage002[75], stage002[76]},
      {stage004[0], stage004[1], stage004[2], stage004[3], stage004[4], stage004[5]},
      {stage006[128], stage005[137], stage004[158], stage003[158], stage002[178]}
   );
   gpc606_5 gpc606_5_97(
      {stage002[77], stage002[78], stage002[79], stage002[80], stage002[81], stage002[82]},
      {stage004[6], stage004[7], stage004[8], stage004[9], stage004[10], stage004[11]},
      {stage006[129], stage005[138], stage004[159], stage003[159], stage002[179]}
   );
   gpc615_5 gpc615_5_98(
      {stage002[83], stage002[84], stage002[85], stage002[86], stage002[87]},
      {stage003[84]},
      {stage004[12], stage004[13], stage004[14], stage004[15], stage004[16], stage004[17]},
      {stage006[130], stage005[139], stage004[160], stage003[160], stage002[180]}
   );
   gpc615_5 gpc615_5_99(
      {stage002[88], stage002[89], stage002[90], stage002[91], stage002[92]},
      {stage003[85]},
      {stage004[18], stage004[19], stage004[20], stage004[21], stage004[22], stage004[23]},
      {stage006[131], stage005[140], stage004[161], stage003[161], stage002[181]}
   );
   gpc615_5 gpc615_5_100(
      {stage002[93], stage002[94], stage002[95], stage002[96], stage002[97]},
      {stage003[86]},
      {stage004[24], stage004[25], stage004[26], stage004[27], stage004[28], stage004[29]},
      {stage006[132], stage005[141], stage004[162], stage003[162], stage002[182]}
   );
   gpc615_5 gpc615_5_101(
      {stage002[98], stage002[99], stage002[100], stage002[101], stage002[102]},
      {stage003[87]},
      {stage004[30], stage004[31], stage004[32], stage004[33], stage004[34], stage004[35]},
      {stage006[133], stage005[142], stage004[163], stage003[163], stage002[183]}
   );
   gpc615_5 gpc615_5_102(
      {stage002[103], stage002[104], stage002[105], stage002[106], stage002[107]},
      {stage003[88]},
      {stage004[36], stage004[37], stage004[38], stage004[39], stage004[40], stage004[41]},
      {stage006[134], stage005[143], stage004[164], stage003[164], stage002[184]}
   );
   gpc615_5 gpc615_5_103(
      {stage002[108], stage002[109], stage002[110], stage002[111], stage002[112]},
      {stage003[89]},
      {stage004[42], stage004[43], stage004[44], stage004[45], stage004[46], stage004[47]},
      {stage006[135], stage005[144], stage004[165], stage003[165], stage002[185]}
   );
   gpc615_5 gpc615_5_104(
      {stage002[113], stage002[114], stage002[115], stage002[116], stage002[117]},
      {stage003[90]},
      {stage004[48], stage004[49], stage004[50], stage004[51], stage004[52], stage004[53]},
      {stage006[136], stage005[145], stage004[166], stage003[166], stage002[186]}
   );
   gpc615_5 gpc615_5_105(
      {stage002[118], stage002[119], stage002[120], stage002[121], stage002[122]},
      {stage003[91]},
      {stage004[54], stage004[55], stage004[56], stage004[57], stage004[58], stage004[59]},
      {stage006[137], stage005[146], stage004[167], stage003[167], stage002[187]}
   );
   gpc615_5 gpc615_5_106(
      {stage002[123], stage002[124], stage002[125], stage002[126], stage002[127]},
      {stage003[92]},
      {stage004[60], stage004[61], stage004[62], stage004[63], stage004[64], stage004[65]},
      {stage006[138], stage005[147], stage004[168], stage003[168], stage002[188]}
   );
   gpc615_5 gpc615_5_107(
      {stage003[93], stage003[94], stage003[95], stage003[96], stage003[97]},
      {stage004[66]},
      {stage005[0], stage005[1], stage005[2], stage005[3], stage005[4], stage005[5]},
      {stage007[128], stage006[139], stage005[148], stage004[169], stage003[169]}
   );
   gpc615_5 gpc615_5_108(
      {stage003[98], stage003[99], stage003[100], stage003[101], stage003[102]},
      {stage004[67]},
      {stage005[6], stage005[7], stage005[8], stage005[9], stage005[10], stage005[11]},
      {stage007[129], stage006[140], stage005[149], stage004[170], stage003[170]}
   );
   gpc615_5 gpc615_5_109(
      {stage003[103], stage003[104], stage003[105], stage003[106], stage003[107]},
      {stage004[68]},
      {stage005[12], stage005[13], stage005[14], stage005[15], stage005[16], stage005[17]},
      {stage007[130], stage006[141], stage005[150], stage004[171], stage003[171]}
   );
   gpc615_5 gpc615_5_110(
      {stage003[108], stage003[109], stage003[110], stage003[111], stage003[112]},
      {stage004[69]},
      {stage005[18], stage005[19], stage005[20], stage005[21], stage005[22], stage005[23]},
      {stage007[131], stage006[142], stage005[151], stage004[172], stage003[172]}
   );
   gpc615_5 gpc615_5_111(
      {stage003[113], stage003[114], stage003[115], stage003[116], stage003[117]},
      {stage004[70]},
      {stage005[24], stage005[25], stage005[26], stage005[27], stage005[28], stage005[29]},
      {stage007[132], stage006[143], stage005[152], stage004[173], stage003[173]}
   );
   gpc615_5 gpc615_5_112(
      {stage003[118], stage003[119], stage003[120], stage003[121], stage003[122]},
      {stage004[71]},
      {stage005[30], stage005[31], stage005[32], stage005[33], stage005[34], stage005[35]},
      {stage007[133], stage006[144], stage005[153], stage004[174], stage003[174]}
   );
   gpc615_5 gpc615_5_113(
      {stage003[123], stage003[124], stage003[125], stage003[126], stage003[127]},
      {stage004[72]},
      {stage005[36], stage005[37], stage005[38], stage005[39], stage005[40], stage005[41]},
      {stage007[134], stage006[145], stage005[154], stage004[175], stage003[175]}
   );
   gpc1_1 gpc1_1_114(
      {stage004[73]},
      {stage004[176]}
   );
   gpc606_5 gpc606_5_115(
      {stage004[74], stage004[75], stage004[76], stage004[77], stage004[78], stage004[79]},
      {stage006[0], stage006[1], stage006[2], stage006[3], stage006[4], stage006[5]},
      {stage008[128], stage007[135], stage006[146], stage005[155], stage004[177]}
   );
   gpc606_5 gpc606_5_116(
      {stage004[80], stage004[81], stage004[82], stage004[83], stage004[84], stage004[85]},
      {stage006[6], stage006[7], stage006[8], stage006[9], stage006[10], stage006[11]},
      {stage008[129], stage007[136], stage006[147], stage005[156], stage004[178]}
   );
   gpc606_5 gpc606_5_117(
      {stage004[86], stage004[87], stage004[88], stage004[89], stage004[90], stage004[91]},
      {stage006[12], stage006[13], stage006[14], stage006[15], stage006[16], stage006[17]},
      {stage008[130], stage007[137], stage006[148], stage005[157], stage004[179]}
   );
   gpc606_5 gpc606_5_118(
      {stage004[92], stage004[93], stage004[94], stage004[95], stage004[96], stage004[97]},
      {stage006[18], stage006[19], stage006[20], stage006[21], stage006[22], stage006[23]},
      {stage008[131], stage007[138], stage006[149], stage005[158], stage004[180]}
   );
   gpc606_5 gpc606_5_119(
      {stage004[98], stage004[99], stage004[100], stage004[101], stage004[102], stage004[103]},
      {stage006[24], stage006[25], stage006[26], stage006[27], stage006[28], stage006[29]},
      {stage008[132], stage007[139], stage006[150], stage005[159], stage004[181]}
   );
   gpc606_5 gpc606_5_120(
      {stage004[104], stage004[105], stage004[106], stage004[107], stage004[108], stage004[109]},
      {stage006[30], stage006[31], stage006[32], stage006[33], stage006[34], stage006[35]},
      {stage008[133], stage007[140], stage006[151], stage005[160], stage004[182]}
   );
   gpc606_5 gpc606_5_121(
      {stage004[110], stage004[111], stage004[112], stage004[113], stage004[114], stage004[115]},
      {stage006[36], stage006[37], stage006[38], stage006[39], stage006[40], stage006[41]},
      {stage008[134], stage007[141], stage006[152], stage005[161], stage004[183]}
   );
   gpc606_5 gpc606_5_122(
      {stage004[116], stage004[117], stage004[118], stage004[119], stage004[120], stage004[121]},
      {stage006[42], stage006[43], stage006[44], stage006[45], stage006[46], stage006[47]},
      {stage008[135], stage007[142], stage006[153], stage005[162], stage004[184]}
   );
   gpc606_5 gpc606_5_123(
      {stage004[122], stage004[123], stage004[124], stage004[125], stage004[126], stage004[127]},
      {stage006[48], stage006[49], stage006[50], stage006[51], stage006[52], stage006[53]},
      {stage008[136], stage007[143], stage006[154], stage005[163], stage004[185]}
   );
   gpc1_1 gpc1_1_124(
      {stage005[42]},
      {stage005[164]}
   );
   gpc1_1 gpc1_1_125(
      {stage005[43]},
      {stage005[165]}
   );
   gpc1_1 gpc1_1_126(
      {stage005[44]},
      {stage005[166]}
   );
   gpc1_1 gpc1_1_127(
      {stage005[45]},
      {stage005[167]}
   );
   gpc1_1 gpc1_1_128(
      {stage005[46]},
      {stage005[168]}
   );
   gpc1_1 gpc1_1_129(
      {stage005[47]},
      {stage005[169]}
   );
   gpc1_1 gpc1_1_130(
      {stage005[48]},
      {stage005[170]}
   );
   gpc1_1 gpc1_1_131(
      {stage005[49]},
      {stage005[171]}
   );
   gpc1_1 gpc1_1_132(
      {stage005[50]},
      {stage005[172]}
   );
   gpc1_1 gpc1_1_133(
      {stage005[51]},
      {stage005[173]}
   );
   gpc1_1 gpc1_1_134(
      {stage005[52]},
      {stage005[174]}
   );
   gpc1_1 gpc1_1_135(
      {stage005[53]},
      {stage005[175]}
   );
   gpc1_1 gpc1_1_136(
      {stage005[54]},
      {stage005[176]}
   );
   gpc1_1 gpc1_1_137(
      {stage005[55]},
      {stage005[177]}
   );
   gpc1_1 gpc1_1_138(
      {stage005[56]},
      {stage005[178]}
   );
   gpc1_1 gpc1_1_139(
      {stage005[57]},
      {stage005[179]}
   );
   gpc1_1 gpc1_1_140(
      {stage005[58]},
      {stage005[180]}
   );
   gpc1_1 gpc1_1_141(
      {stage005[59]},
      {stage005[181]}
   );
   gpc1_1 gpc1_1_142(
      {stage005[60]},
      {stage005[182]}
   );
   gpc1_1 gpc1_1_143(
      {stage005[61]},
      {stage005[183]}
   );
   gpc1_1 gpc1_1_144(
      {stage005[62]},
      {stage005[184]}
   );
   gpc1_1 gpc1_1_145(
      {stage005[63]},
      {stage005[185]}
   );
   gpc1_1 gpc1_1_146(
      {stage005[64]},
      {stage005[186]}
   );
   gpc1_1 gpc1_1_147(
      {stage005[65]},
      {stage005[187]}
   );
   gpc1_1 gpc1_1_148(
      {stage005[66]},
      {stage005[188]}
   );
   gpc1_1 gpc1_1_149(
      {stage005[67]},
      {stage005[189]}
   );
   gpc1_1 gpc1_1_150(
      {stage005[68]},
      {stage005[190]}
   );
   gpc1_1 gpc1_1_151(
      {stage005[69]},
      {stage005[191]}
   );
   gpc1_1 gpc1_1_152(
      {stage005[70]},
      {stage005[192]}
   );
   gpc1_1 gpc1_1_153(
      {stage005[71]},
      {stage005[193]}
   );
   gpc1_1 gpc1_1_154(
      {stage005[72]},
      {stage005[194]}
   );
   gpc1_1 gpc1_1_155(
      {stage005[73]},
      {stage005[195]}
   );
   gpc1_1 gpc1_1_156(
      {stage005[74]},
      {stage005[196]}
   );
   gpc1_1 gpc1_1_157(
      {stage005[75]},
      {stage005[197]}
   );
   gpc1_1 gpc1_1_158(
      {stage005[76]},
      {stage005[198]}
   );
   gpc1_1 gpc1_1_159(
      {stage005[77]},
      {stage005[199]}
   );
   gpc1_1 gpc1_1_160(
      {stage005[78]},
      {stage005[200]}
   );
   gpc1_1 gpc1_1_161(
      {stage005[79]},
      {stage005[201]}
   );
   gpc1_1 gpc1_1_162(
      {stage005[80]},
      {stage005[202]}
   );
   gpc1_1 gpc1_1_163(
      {stage005[81]},
      {stage005[203]}
   );
   gpc606_5 gpc606_5_164(
      {stage005[82], stage005[83], stage005[84], stage005[85], stage005[86], stage005[87]},
      {stage007[0], stage007[1], stage007[2], stage007[3], stage007[4], stage007[5]},
      {stage009[128], stage008[137], stage007[144], stage006[155], stage005[204]}
   );
   gpc615_5 gpc615_5_165(
      {stage005[88], stage005[89], stage005[90], stage005[91], stage005[92]},
      {stage006[54]},
      {stage007[6], stage007[7], stage007[8], stage007[9], stage007[10], stage007[11]},
      {stage009[129], stage008[138], stage007[145], stage006[156], stage005[205]}
   );
   gpc615_5 gpc615_5_166(
      {stage005[93], stage005[94], stage005[95], stage005[96], stage005[97]},
      {stage006[55]},
      {stage007[12], stage007[13], stage007[14], stage007[15], stage007[16], stage007[17]},
      {stage009[130], stage008[139], stage007[146], stage006[157], stage005[206]}
   );
   gpc615_5 gpc615_5_167(
      {stage005[98], stage005[99], stage005[100], stage005[101], stage005[102]},
      {stage006[56]},
      {stage007[18], stage007[19], stage007[20], stage007[21], stage007[22], stage007[23]},
      {stage009[131], stage008[140], stage007[147], stage006[158], stage005[207]}
   );
   gpc615_5 gpc615_5_168(
      {stage005[103], stage005[104], stage005[105], stage005[106], stage005[107]},
      {stage006[57]},
      {stage007[24], stage007[25], stage007[26], stage007[27], stage007[28], stage007[29]},
      {stage009[132], stage008[141], stage007[148], stage006[159], stage005[208]}
   );
   gpc615_5 gpc615_5_169(
      {stage005[108], stage005[109], stage005[110], stage005[111], stage005[112]},
      {stage006[58]},
      {stage007[30], stage007[31], stage007[32], stage007[33], stage007[34], stage007[35]},
      {stage009[133], stage008[142], stage007[149], stage006[160], stage005[209]}
   );
   gpc615_5 gpc615_5_170(
      {stage005[113], stage005[114], stage005[115], stage005[116], stage005[117]},
      {stage006[59]},
      {stage007[36], stage007[37], stage007[38], stage007[39], stage007[40], stage007[41]},
      {stage009[134], stage008[143], stage007[150], stage006[161], stage005[210]}
   );
   gpc615_5 gpc615_5_171(
      {stage005[118], stage005[119], stage005[120], stage005[121], stage005[122]},
      {stage006[60]},
      {stage007[42], stage007[43], stage007[44], stage007[45], stage007[46], stage007[47]},
      {stage009[135], stage008[144], stage007[151], stage006[162], stage005[211]}
   );
   gpc615_5 gpc615_5_172(
      {stage005[123], stage005[124], stage005[125], stage005[126], stage005[127]},
      {stage006[61]},
      {stage007[48], stage007[49], stage007[50], stage007[51], stage007[52], stage007[53]},
      {stage009[136], stage008[145], stage007[152], stage006[163], stage005[212]}
   );
   gpc1_1 gpc1_1_173(
      {stage006[62]},
      {stage006[164]}
   );
   gpc1_1 gpc1_1_174(
      {stage006[63]},
      {stage006[165]}
   );
   gpc1_1 gpc1_1_175(
      {stage006[64]},
      {stage006[166]}
   );
   gpc1_1 gpc1_1_176(
      {stage006[65]},
      {stage006[167]}
   );
   gpc1_1 gpc1_1_177(
      {stage006[66]},
      {stage006[168]}
   );
   gpc1_1 gpc1_1_178(
      {stage006[67]},
      {stage006[169]}
   );
   gpc1_1 gpc1_1_179(
      {stage006[68]},
      {stage006[170]}
   );
   gpc1_1 gpc1_1_180(
      {stage006[69]},
      {stage006[171]}
   );
   gpc1_1 gpc1_1_181(
      {stage006[70]},
      {stage006[172]}
   );
   gpc1_1 gpc1_1_182(
      {stage006[71]},
      {stage006[173]}
   );
   gpc1_1 gpc1_1_183(
      {stage006[72]},
      {stage006[174]}
   );
   gpc1_1 gpc1_1_184(
      {stage006[73]},
      {stage006[175]}
   );
   gpc1_1 gpc1_1_185(
      {stage006[74]},
      {stage006[176]}
   );
   gpc1_1 gpc1_1_186(
      {stage006[75]},
      {stage006[177]}
   );
   gpc606_5 gpc606_5_187(
      {stage006[76], stage006[77], stage006[78], stage006[79], stage006[80], stage006[81]},
      {stage008[0], stage008[1], stage008[2], stage008[3], stage008[4], stage008[5]},
      {stage010[128], stage009[137], stage008[146], stage007[153], stage006[178]}
   );
   gpc606_5 gpc606_5_188(
      {stage006[82], stage006[83], stage006[84], stage006[85], stage006[86], stage006[87]},
      {stage008[6], stage008[7], stage008[8], stage008[9], stage008[10], stage008[11]},
      {stage010[129], stage009[138], stage008[147], stage007[154], stage006[179]}
   );
   gpc615_5 gpc615_5_189(
      {stage006[88], stage006[89], stage006[90], stage006[91], stage006[92]},
      {stage007[54]},
      {stage008[12], stage008[13], stage008[14], stage008[15], stage008[16], stage008[17]},
      {stage010[130], stage009[139], stage008[148], stage007[155], stage006[180]}
   );
   gpc615_5 gpc615_5_190(
      {stage006[93], stage006[94], stage006[95], stage006[96], stage006[97]},
      {stage007[55]},
      {stage008[18], stage008[19], stage008[20], stage008[21], stage008[22], stage008[23]},
      {stage010[131], stage009[140], stage008[149], stage007[156], stage006[181]}
   );
   gpc615_5 gpc615_5_191(
      {stage006[98], stage006[99], stage006[100], stage006[101], stage006[102]},
      {stage007[56]},
      {stage008[24], stage008[25], stage008[26], stage008[27], stage008[28], stage008[29]},
      {stage010[132], stage009[141], stage008[150], stage007[157], stage006[182]}
   );
   gpc615_5 gpc615_5_192(
      {stage006[103], stage006[104], stage006[105], stage006[106], stage006[107]},
      {stage007[57]},
      {stage008[30], stage008[31], stage008[32], stage008[33], stage008[34], stage008[35]},
      {stage010[133], stage009[142], stage008[151], stage007[158], stage006[183]}
   );
   gpc615_5 gpc615_5_193(
      {stage006[108], stage006[109], stage006[110], stage006[111], stage006[112]},
      {stage007[58]},
      {stage008[36], stage008[37], stage008[38], stage008[39], stage008[40], stage008[41]},
      {stage010[134], stage009[143], stage008[152], stage007[159], stage006[184]}
   );
   gpc615_5 gpc615_5_194(
      {stage006[113], stage006[114], stage006[115], stage006[116], stage006[117]},
      {stage007[59]},
      {stage008[42], stage008[43], stage008[44], stage008[45], stage008[46], stage008[47]},
      {stage010[135], stage009[144], stage008[153], stage007[160], stage006[185]}
   );
   gpc615_5 gpc615_5_195(
      {stage006[118], stage006[119], stage006[120], stage006[121], stage006[122]},
      {stage007[60]},
      {stage008[48], stage008[49], stage008[50], stage008[51], stage008[52], stage008[53]},
      {stage010[136], stage009[145], stage008[154], stage007[161], stage006[186]}
   );
   gpc615_5 gpc615_5_196(
      {stage006[123], stage006[124], stage006[125], stage006[126], stage006[127]},
      {stage007[61]},
      {stage008[54], stage008[55], stage008[56], stage008[57], stage008[58], stage008[59]},
      {stage010[137], stage009[146], stage008[155], stage007[162], stage006[187]}
   );
   gpc1_1 gpc1_1_197(
      {stage007[62]},
      {stage007[163]}
   );
   gpc1_1 gpc1_1_198(
      {stage007[63]},
      {stage007[164]}
   );
   gpc1_1 gpc1_1_199(
      {stage007[64]},
      {stage007[165]}
   );
   gpc1_1 gpc1_1_200(
      {stage007[65]},
      {stage007[166]}
   );
   gpc1_1 gpc1_1_201(
      {stage007[66]},
      {stage007[167]}
   );
   gpc1_1 gpc1_1_202(
      {stage007[67]},
      {stage007[168]}
   );
   gpc1_1 gpc1_1_203(
      {stage007[68]},
      {stage007[169]}
   );
   gpc1_1 gpc1_1_204(
      {stage007[69]},
      {stage007[170]}
   );
   gpc1_1 gpc1_1_205(
      {stage007[70]},
      {stage007[171]}
   );
   gpc1_1 gpc1_1_206(
      {stage007[71]},
      {stage007[172]}
   );
   gpc1_1 gpc1_1_207(
      {stage007[72]},
      {stage007[173]}
   );
   gpc1_1 gpc1_1_208(
      {stage007[73]},
      {stage007[174]}
   );
   gpc1_1 gpc1_1_209(
      {stage007[74]},
      {stage007[175]}
   );
   gpc1_1 gpc1_1_210(
      {stage007[75]},
      {stage007[176]}
   );
   gpc1_1 gpc1_1_211(
      {stage007[76]},
      {stage007[177]}
   );
   gpc1_1 gpc1_1_212(
      {stage007[77]},
      {stage007[178]}
   );
   gpc1_1 gpc1_1_213(
      {stage007[78]},
      {stage007[179]}
   );
   gpc1_1 gpc1_1_214(
      {stage007[79]},
      {stage007[180]}
   );
   gpc1_1 gpc1_1_215(
      {stage007[80]},
      {stage007[181]}
   );
   gpc1_1 gpc1_1_216(
      {stage007[81]},
      {stage007[182]}
   );
   gpc1_1 gpc1_1_217(
      {stage007[82]},
      {stage007[183]}
   );
   gpc615_5 gpc615_5_218(
      {stage007[83], stage007[84], stage007[85], stage007[86], stage007[87]},
      {stage008[60]},
      {stage009[0], stage009[1], stage009[2], stage009[3], stage009[4], stage009[5]},
      {stage011[128], stage010[138], stage009[147], stage008[156], stage007[184]}
   );
   gpc615_5 gpc615_5_219(
      {stage007[88], stage007[89], stage007[90], stage007[91], stage007[92]},
      {stage008[61]},
      {stage009[6], stage009[7], stage009[8], stage009[9], stage009[10], stage009[11]},
      {stage011[129], stage010[139], stage009[148], stage008[157], stage007[185]}
   );
   gpc615_5 gpc615_5_220(
      {stage007[93], stage007[94], stage007[95], stage007[96], stage007[97]},
      {stage008[62]},
      {stage009[12], stage009[13], stage009[14], stage009[15], stage009[16], stage009[17]},
      {stage011[130], stage010[140], stage009[149], stage008[158], stage007[186]}
   );
   gpc615_5 gpc615_5_221(
      {stage007[98], stage007[99], stage007[100], stage007[101], stage007[102]},
      {stage008[63]},
      {stage009[18], stage009[19], stage009[20], stage009[21], stage009[22], stage009[23]},
      {stage011[131], stage010[141], stage009[150], stage008[159], stage007[187]}
   );
   gpc615_5 gpc615_5_222(
      {stage007[103], stage007[104], stage007[105], stage007[106], stage007[107]},
      {stage008[64]},
      {stage009[24], stage009[25], stage009[26], stage009[27], stage009[28], stage009[29]},
      {stage011[132], stage010[142], stage009[151], stage008[160], stage007[188]}
   );
   gpc615_5 gpc615_5_223(
      {stage007[108], stage007[109], stage007[110], stage007[111], stage007[112]},
      {stage008[65]},
      {stage009[30], stage009[31], stage009[32], stage009[33], stage009[34], stage009[35]},
      {stage011[133], stage010[143], stage009[152], stage008[161], stage007[189]}
   );
   gpc615_5 gpc615_5_224(
      {stage007[113], stage007[114], stage007[115], stage007[116], stage007[117]},
      {stage008[66]},
      {stage009[36], stage009[37], stage009[38], stage009[39], stage009[40], stage009[41]},
      {stage011[134], stage010[144], stage009[153], stage008[162], stage007[190]}
   );
   gpc615_5 gpc615_5_225(
      {stage007[118], stage007[119], stage007[120], stage007[121], stage007[122]},
      {stage008[67]},
      {stage009[42], stage009[43], stage009[44], stage009[45], stage009[46], stage009[47]},
      {stage011[135], stage010[145], stage009[154], stage008[163], stage007[191]}
   );
   gpc615_5 gpc615_5_226(
      {stage007[123], stage007[124], stage007[125], stage007[126], stage007[127]},
      {stage008[68]},
      {stage009[48], stage009[49], stage009[50], stage009[51], stage009[52], stage009[53]},
      {stage011[136], stage010[146], stage009[155], stage008[164], stage007[192]}
   );
   gpc606_5 gpc606_5_227(
      {stage008[69], stage008[70], stage008[71], stage008[72], stage008[73], stage008[74]},
      {stage010[0], stage010[1], stage010[2], stage010[3], stage010[4], stage010[5]},
      {stage012[128], stage011[137], stage010[147], stage009[156], stage008[165]}
   );
   gpc606_5 gpc606_5_228(
      {stage008[75], stage008[76], stage008[77], stage008[78], stage008[79], stage008[80]},
      {stage010[6], stage010[7], stage010[8], stage010[9], stage010[10], stage010[11]},
      {stage012[129], stage011[138], stage010[148], stage009[157], stage008[166]}
   );
   gpc606_5 gpc606_5_229(
      {stage008[81], stage008[82], stage008[83], stage008[84], stage008[85], stage008[86]},
      {stage010[12], stage010[13], stage010[14], stage010[15], stage010[16], stage010[17]},
      {stage012[130], stage011[139], stage010[149], stage009[158], stage008[167]}
   );
   gpc606_5 gpc606_5_230(
      {stage008[87], stage008[88], stage008[89], stage008[90], stage008[91], stage008[92]},
      {stage010[18], stage010[19], stage010[20], stage010[21], stage010[22], stage010[23]},
      {stage012[131], stage011[140], stage010[150], stage009[159], stage008[168]}
   );
   gpc615_5 gpc615_5_231(
      {stage008[93], stage008[94], stage008[95], stage008[96], stage008[97]},
      {stage009[54]},
      {stage010[24], stage010[25], stage010[26], stage010[27], stage010[28], stage010[29]},
      {stage012[132], stage011[141], stage010[151], stage009[160], stage008[169]}
   );
   gpc615_5 gpc615_5_232(
      {stage008[98], stage008[99], stage008[100], stage008[101], stage008[102]},
      {stage009[55]},
      {stage010[30], stage010[31], stage010[32], stage010[33], stage010[34], stage010[35]},
      {stage012[133], stage011[142], stage010[152], stage009[161], stage008[170]}
   );
   gpc615_5 gpc615_5_233(
      {stage008[103], stage008[104], stage008[105], stage008[106], stage008[107]},
      {stage009[56]},
      {stage010[36], stage010[37], stage010[38], stage010[39], stage010[40], stage010[41]},
      {stage012[134], stage011[143], stage010[153], stage009[162], stage008[171]}
   );
   gpc615_5 gpc615_5_234(
      {stage008[108], stage008[109], stage008[110], stage008[111], stage008[112]},
      {stage009[57]},
      {stage010[42], stage010[43], stage010[44], stage010[45], stage010[46], stage010[47]},
      {stage012[135], stage011[144], stage010[154], stage009[163], stage008[172]}
   );
   gpc615_5 gpc615_5_235(
      {stage008[113], stage008[114], stage008[115], stage008[116], stage008[117]},
      {stage009[58]},
      {stage010[48], stage010[49], stage010[50], stage010[51], stage010[52], stage010[53]},
      {stage012[136], stage011[145], stage010[155], stage009[164], stage008[173]}
   );
   gpc615_5 gpc615_5_236(
      {stage008[118], stage008[119], stage008[120], stage008[121], stage008[122]},
      {stage009[59]},
      {stage010[54], stage010[55], stage010[56], stage010[57], stage010[58], stage010[59]},
      {stage012[137], stage011[146], stage010[156], stage009[165], stage008[174]}
   );
   gpc615_5 gpc615_5_237(
      {stage008[123], stage008[124], stage008[125], stage008[126], stage008[127]},
      {stage009[60]},
      {stage010[60], stage010[61], stage010[62], stage010[63], stage010[64], stage010[65]},
      {stage012[138], stage011[147], stage010[157], stage009[166], stage008[175]}
   );
   gpc1_1 gpc1_1_238(
      {stage009[61]},
      {stage009[167]}
   );
   gpc1_1 gpc1_1_239(
      {stage009[62]},
      {stage009[168]}
   );
   gpc1_1 gpc1_1_240(
      {stage009[63]},
      {stage009[169]}
   );
   gpc1_1 gpc1_1_241(
      {stage009[64]},
      {stage009[170]}
   );
   gpc1_1 gpc1_1_242(
      {stage009[65]},
      {stage009[171]}
   );
   gpc1_1 gpc1_1_243(
      {stage009[66]},
      {stage009[172]}
   );
   gpc1_1 gpc1_1_244(
      {stage009[67]},
      {stage009[173]}
   );
   gpc1_1 gpc1_1_245(
      {stage009[68]},
      {stage009[174]}
   );
   gpc1_1 gpc1_1_246(
      {stage009[69]},
      {stage009[175]}
   );
   gpc1_1 gpc1_1_247(
      {stage009[70]},
      {stage009[176]}
   );
   gpc606_5 gpc606_5_248(
      {stage009[71], stage009[72], stage009[73], stage009[74], stage009[75], stage009[76]},
      {stage011[0], stage011[1], stage011[2], stage011[3], stage011[4], stage011[5]},
      {stage013[128], stage012[139], stage011[148], stage010[158], stage009[177]}
   );
   gpc606_5 gpc606_5_249(
      {stage009[77], stage009[78], stage009[79], stage009[80], stage009[81], stage009[82]},
      {stage011[6], stage011[7], stage011[8], stage011[9], stage011[10], stage011[11]},
      {stage013[129], stage012[140], stage011[149], stage010[159], stage009[178]}
   );
   gpc615_5 gpc615_5_250(
      {stage009[83], stage009[84], stage009[85], stage009[86], stage009[87]},
      {stage010[66]},
      {stage011[12], stage011[13], stage011[14], stage011[15], stage011[16], stage011[17]},
      {stage013[130], stage012[141], stage011[150], stage010[160], stage009[179]}
   );
   gpc615_5 gpc615_5_251(
      {stage009[88], stage009[89], stage009[90], stage009[91], stage009[92]},
      {stage010[67]},
      {stage011[18], stage011[19], stage011[20], stage011[21], stage011[22], stage011[23]},
      {stage013[131], stage012[142], stage011[151], stage010[161], stage009[180]}
   );
   gpc615_5 gpc615_5_252(
      {stage009[93], stage009[94], stage009[95], stage009[96], stage009[97]},
      {stage010[68]},
      {stage011[24], stage011[25], stage011[26], stage011[27], stage011[28], stage011[29]},
      {stage013[132], stage012[143], stage011[152], stage010[162], stage009[181]}
   );
   gpc615_5 gpc615_5_253(
      {stage009[98], stage009[99], stage009[100], stage009[101], stage009[102]},
      {stage010[69]},
      {stage011[30], stage011[31], stage011[32], stage011[33], stage011[34], stage011[35]},
      {stage013[133], stage012[144], stage011[153], stage010[163], stage009[182]}
   );
   gpc615_5 gpc615_5_254(
      {stage009[103], stage009[104], stage009[105], stage009[106], stage009[107]},
      {stage010[70]},
      {stage011[36], stage011[37], stage011[38], stage011[39], stage011[40], stage011[41]},
      {stage013[134], stage012[145], stage011[154], stage010[164], stage009[183]}
   );
   gpc615_5 gpc615_5_255(
      {stage009[108], stage009[109], stage009[110], stage009[111], stage009[112]},
      {stage010[71]},
      {stage011[42], stage011[43], stage011[44], stage011[45], stage011[46], stage011[47]},
      {stage013[135], stage012[146], stage011[155], stage010[165], stage009[184]}
   );
   gpc615_5 gpc615_5_256(
      {stage009[113], stage009[114], stage009[115], stage009[116], stage009[117]},
      {stage010[72]},
      {stage011[48], stage011[49], stage011[50], stage011[51], stage011[52], stage011[53]},
      {stage013[136], stage012[147], stage011[156], stage010[166], stage009[185]}
   );
   gpc615_5 gpc615_5_257(
      {stage009[118], stage009[119], stage009[120], stage009[121], stage009[122]},
      {stage010[73]},
      {stage011[54], stage011[55], stage011[56], stage011[57], stage011[58], stage011[59]},
      {stage013[137], stage012[148], stage011[157], stage010[167], stage009[186]}
   );
   gpc615_5 gpc615_5_258(
      {stage009[123], stage009[124], stage009[125], stage009[126], stage009[127]},
      {stage010[74]},
      {stage011[60], stage011[61], stage011[62], stage011[63], stage011[64], stage011[65]},
      {stage013[138], stage012[149], stage011[158], stage010[168], stage009[187]}
   );
   gpc1_1 gpc1_1_259(
      {stage010[75]},
      {stage010[169]}
   );
   gpc1_1 gpc1_1_260(
      {stage010[76]},
      {stage010[170]}
   );
   gpc1_1 gpc1_1_261(
      {stage010[77]},
      {stage010[171]}
   );
   gpc1_1 gpc1_1_262(
      {stage010[78]},
      {stage010[172]}
   );
   gpc1_1 gpc1_1_263(
      {stage010[79]},
      {stage010[173]}
   );
   gpc1_1 gpc1_1_264(
      {stage010[80]},
      {stage010[174]}
   );
   gpc1_1 gpc1_1_265(
      {stage010[81]},
      {stage010[175]}
   );
   gpc1_1 gpc1_1_266(
      {stage010[82]},
      {stage010[176]}
   );
   gpc1_1 gpc1_1_267(
      {stage010[83]},
      {stage010[177]}
   );
   gpc1_1 gpc1_1_268(
      {stage010[84]},
      {stage010[178]}
   );
   gpc1_1 gpc1_1_269(
      {stage010[85]},
      {stage010[179]}
   );
   gpc1_1 gpc1_1_270(
      {stage010[86]},
      {stage010[180]}
   );
   gpc606_5 gpc606_5_271(
      {stage010[87], stage010[88], stage010[89], stage010[90], stage010[91], stage010[92]},
      {stage012[0], stage012[1], stage012[2], stage012[3], stage012[4], stage012[5]},
      {stage014[128], stage013[139], stage012[150], stage011[159], stage010[181]}
   );
   gpc606_5 gpc606_5_272(
      {stage010[93], stage010[94], stage010[95], stage010[96], stage010[97], stage010[98]},
      {stage012[6], stage012[7], stage012[8], stage012[9], stage012[10], stage012[11]},
      {stage014[129], stage013[140], stage012[151], stage011[160], stage010[182]}
   );
   gpc606_5 gpc606_5_273(
      {stage010[99], stage010[100], stage010[101], stage010[102], stage010[103], stage010[104]},
      {stage012[12], stage012[13], stage012[14], stage012[15], stage012[16], stage012[17]},
      {stage014[130], stage013[141], stage012[152], stage011[161], stage010[183]}
   );
   gpc606_5 gpc606_5_274(
      {stage010[105], stage010[106], stage010[107], stage010[108], stage010[109], stage010[110]},
      {stage012[18], stage012[19], stage012[20], stage012[21], stage012[22], stage012[23]},
      {stage014[131], stage013[142], stage012[153], stage011[162], stage010[184]}
   );
   gpc606_5 gpc606_5_275(
      {stage010[111], stage010[112], stage010[113], stage010[114], stage010[115], stage010[116]},
      {stage012[24], stage012[25], stage012[26], stage012[27], stage012[28], stage012[29]},
      {stage014[132], stage013[143], stage012[154], stage011[163], stage010[185]}
   );
   gpc606_5 gpc606_5_276(
      {stage010[117], stage010[118], stage010[119], stage010[120], stage010[121], stage010[122]},
      {stage012[30], stage012[31], stage012[32], stage012[33], stage012[34], stage012[35]},
      {stage014[133], stage013[144], stage012[155], stage011[164], stage010[186]}
   );
   gpc615_5 gpc615_5_277(
      {stage010[123], stage010[124], stage010[125], stage010[126], stage010[127]},
      {stage011[66]},
      {stage012[36], stage012[37], stage012[38], stage012[39], stage012[40], stage012[41]},
      {stage014[134], stage013[145], stage012[156], stage011[165], stage010[187]}
   );
   gpc1_1 gpc1_1_278(
      {stage011[67]},
      {stage011[166]}
   );
   gpc1_1 gpc1_1_279(
      {stage011[68]},
      {stage011[167]}
   );
   gpc1_1 gpc1_1_280(
      {stage011[69]},
      {stage011[168]}
   );
   gpc1_1 gpc1_1_281(
      {stage011[70]},
      {stage011[169]}
   );
   gpc1_1 gpc1_1_282(
      {stage011[71]},
      {stage011[170]}
   );
   gpc1_1 gpc1_1_283(
      {stage011[72]},
      {stage011[171]}
   );
   gpc1_1 gpc1_1_284(
      {stage011[73]},
      {stage011[172]}
   );
   gpc1_1 gpc1_1_285(
      {stage011[74]},
      {stage011[173]}
   );
   gpc1_1 gpc1_1_286(
      {stage011[75]},
      {stage011[174]}
   );
   gpc1_1 gpc1_1_287(
      {stage011[76]},
      {stage011[175]}
   );
   gpc1_1 gpc1_1_288(
      {stage011[77]},
      {stage011[176]}
   );
   gpc1_1 gpc1_1_289(
      {stage011[78]},
      {stage011[177]}
   );
   gpc1_1 gpc1_1_290(
      {stage011[79]},
      {stage011[178]}
   );
   gpc1_1 gpc1_1_291(
      {stage011[80]},
      {stage011[179]}
   );
   gpc1_1 gpc1_1_292(
      {stage011[81]},
      {stage011[180]}
   );
   gpc1_1 gpc1_1_293(
      {stage011[82]},
      {stage011[181]}
   );
   gpc1_1 gpc1_1_294(
      {stage011[83]},
      {stage011[182]}
   );
   gpc1_1 gpc1_1_295(
      {stage011[84]},
      {stage011[183]}
   );
   gpc1_1 gpc1_1_296(
      {stage011[85]},
      {stage011[184]}
   );
   gpc1_1 gpc1_1_297(
      {stage011[86]},
      {stage011[185]}
   );
   gpc1_1 gpc1_1_298(
      {stage011[87]},
      {stage011[186]}
   );
   gpc1_1 gpc1_1_299(
      {stage011[88]},
      {stage011[187]}
   );
   gpc1_1 gpc1_1_300(
      {stage011[89]},
      {stage011[188]}
   );
   gpc1_1 gpc1_1_301(
      {stage011[90]},
      {stage011[189]}
   );
   gpc1_1 gpc1_1_302(
      {stage011[91]},
      {stage011[190]}
   );
   gpc1_1 gpc1_1_303(
      {stage011[92]},
      {stage011[191]}
   );
   gpc1_1 gpc1_1_304(
      {stage011[93]},
      {stage011[192]}
   );
   gpc1_1 gpc1_1_305(
      {stage011[94]},
      {stage011[193]}
   );
   gpc1_1 gpc1_1_306(
      {stage011[95]},
      {stage011[194]}
   );
   gpc1_1 gpc1_1_307(
      {stage011[96]},
      {stage011[195]}
   );
   gpc606_5 gpc606_5_308(
      {stage011[97], stage011[98], stage011[99], stage011[100], stage011[101], stage011[102]},
      {stage013[0], stage013[1], stage013[2], stage013[3], stage013[4], stage013[5]},
      {stage015[128], stage014[135], stage013[146], stage012[157], stage011[196]}
   );
   gpc615_5 gpc615_5_309(
      {stage011[103], stage011[104], stage011[105], stage011[106], stage011[107]},
      {stage012[42]},
      {stage013[6], stage013[7], stage013[8], stage013[9], stage013[10], stage013[11]},
      {stage015[129], stage014[136], stage013[147], stage012[158], stage011[197]}
   );
   gpc615_5 gpc615_5_310(
      {stage011[108], stage011[109], stage011[110], stage011[111], stage011[112]},
      {stage012[43]},
      {stage013[12], stage013[13], stage013[14], stage013[15], stage013[16], stage013[17]},
      {stage015[130], stage014[137], stage013[148], stage012[159], stage011[198]}
   );
   gpc615_5 gpc615_5_311(
      {stage011[113], stage011[114], stage011[115], stage011[116], stage011[117]},
      {stage012[44]},
      {stage013[18], stage013[19], stage013[20], stage013[21], stage013[22], stage013[23]},
      {stage015[131], stage014[138], stage013[149], stage012[160], stage011[199]}
   );
   gpc615_5 gpc615_5_312(
      {stage011[118], stage011[119], stage011[120], stage011[121], stage011[122]},
      {stage012[45]},
      {stage013[24], stage013[25], stage013[26], stage013[27], stage013[28], stage013[29]},
      {stage015[132], stage014[139], stage013[150], stage012[161], stage011[200]}
   );
   gpc615_5 gpc615_5_313(
      {stage011[123], stage011[124], stage011[125], stage011[126], stage011[127]},
      {stage012[46]},
      {stage013[30], stage013[31], stage013[32], stage013[33], stage013[34], stage013[35]},
      {stage015[133], stage014[140], stage013[151], stage012[162], stage011[201]}
   );
   gpc1_1 gpc1_1_314(
      {stage012[47]},
      {stage012[163]}
   );
   gpc1_1 gpc1_1_315(
      {stage012[48]},
      {stage012[164]}
   );
   gpc1_1 gpc1_1_316(
      {stage012[49]},
      {stage012[165]}
   );
   gpc1_1 gpc1_1_317(
      {stage012[50]},
      {stage012[166]}
   );
   gpc1_1 gpc1_1_318(
      {stage012[51]},
      {stage012[167]}
   );
   gpc1_1 gpc1_1_319(
      {stage012[52]},
      {stage012[168]}
   );
   gpc1_1 gpc1_1_320(
      {stage012[53]},
      {stage012[169]}
   );
   gpc1_1 gpc1_1_321(
      {stage012[54]},
      {stage012[170]}
   );
   gpc1_1 gpc1_1_322(
      {stage012[55]},
      {stage012[171]}
   );
   gpc1_1 gpc1_1_323(
      {stage012[56]},
      {stage012[172]}
   );
   gpc1_1 gpc1_1_324(
      {stage012[57]},
      {stage012[173]}
   );
   gpc1_1 gpc1_1_325(
      {stage012[58]},
      {stage012[174]}
   );
   gpc1_1 gpc1_1_326(
      {stage012[59]},
      {stage012[175]}
   );
   gpc1_1 gpc1_1_327(
      {stage012[60]},
      {stage012[176]}
   );
   gpc1_1 gpc1_1_328(
      {stage012[61]},
      {stage012[177]}
   );
   gpc1_1 gpc1_1_329(
      {stage012[62]},
      {stage012[178]}
   );
   gpc1_1 gpc1_1_330(
      {stage012[63]},
      {stage012[179]}
   );
   gpc1_1 gpc1_1_331(
      {stage012[64]},
      {stage012[180]}
   );
   gpc1_1 gpc1_1_332(
      {stage012[65]},
      {stage012[181]}
   );
   gpc1_1 gpc1_1_333(
      {stage012[66]},
      {stage012[182]}
   );
   gpc1_1 gpc1_1_334(
      {stage012[67]},
      {stage012[183]}
   );
   gpc1_1 gpc1_1_335(
      {stage012[68]},
      {stage012[184]}
   );
   gpc1_1 gpc1_1_336(
      {stage012[69]},
      {stage012[185]}
   );
   gpc1_1 gpc1_1_337(
      {stage012[70]},
      {stage012[186]}
   );
   gpc1_1 gpc1_1_338(
      {stage012[71]},
      {stage012[187]}
   );
   gpc1_1 gpc1_1_339(
      {stage012[72]},
      {stage012[188]}
   );
   gpc1_1 gpc1_1_340(
      {stage012[73]},
      {stage012[189]}
   );
   gpc1_1 gpc1_1_341(
      {stage012[74]},
      {stage012[190]}
   );
   gpc1_1 gpc1_1_342(
      {stage012[75]},
      {stage012[191]}
   );
   gpc1_1 gpc1_1_343(
      {stage012[76]},
      {stage012[192]}
   );
   gpc1_1 gpc1_1_344(
      {stage012[77]},
      {stage012[193]}
   );
   gpc1_1 gpc1_1_345(
      {stage012[78]},
      {stage012[194]}
   );
   gpc1_1 gpc1_1_346(
      {stage012[79]},
      {stage012[195]}
   );
   gpc1_1 gpc1_1_347(
      {stage012[80]},
      {stage012[196]}
   );
   gpc1_1 gpc1_1_348(
      {stage012[81]},
      {stage012[197]}
   );
   gpc1_1 gpc1_1_349(
      {stage012[82]},
      {stage012[198]}
   );
   gpc1_1 gpc1_1_350(
      {stage012[83]},
      {stage012[199]}
   );
   gpc1_1 gpc1_1_351(
      {stage012[84]},
      {stage012[200]}
   );
   gpc1_1 gpc1_1_352(
      {stage012[85]},
      {stage012[201]}
   );
   gpc1_1 gpc1_1_353(
      {stage012[86]},
      {stage012[202]}
   );
   gpc1_1 gpc1_1_354(
      {stage012[87]},
      {stage012[203]}
   );
   gpc1_1 gpc1_1_355(
      {stage012[88]},
      {stage012[204]}
   );
   gpc1_1 gpc1_1_356(
      {stage012[89]},
      {stage012[205]}
   );
   gpc1_1 gpc1_1_357(
      {stage012[90]},
      {stage012[206]}
   );
   gpc1_1 gpc1_1_358(
      {stage012[91]},
      {stage012[207]}
   );
   gpc1_1 gpc1_1_359(
      {stage012[92]},
      {stage012[208]}
   );
   gpc1_1 gpc1_1_360(
      {stage012[93]},
      {stage012[209]}
   );
   gpc1_1 gpc1_1_361(
      {stage012[94]},
      {stage012[210]}
   );
   gpc1_1 gpc1_1_362(
      {stage012[95]},
      {stage012[211]}
   );
   gpc1_1 gpc1_1_363(
      {stage012[96]},
      {stage012[212]}
   );
   gpc1_1 gpc1_1_364(
      {stage012[97]},
      {stage012[213]}
   );
   gpc615_5 gpc615_5_365(
      {stage012[98], stage012[99], stage012[100], stage012[101], stage012[102]},
      {stage013[36]},
      {stage014[0], stage014[1], stage014[2], stage014[3], stage014[4], stage014[5]},
      {stage016[128], stage015[134], stage014[141], stage013[152], stage012[214]}
   );
   gpc615_5 gpc615_5_366(
      {stage012[103], stage012[104], stage012[105], stage012[106], stage012[107]},
      {stage013[37]},
      {stage014[6], stage014[7], stage014[8], stage014[9], stage014[10], stage014[11]},
      {stage016[129], stage015[135], stage014[142], stage013[153], stage012[215]}
   );
   gpc615_5 gpc615_5_367(
      {stage012[108], stage012[109], stage012[110], stage012[111], stage012[112]},
      {stage013[38]},
      {stage014[12], stage014[13], stage014[14], stage014[15], stage014[16], stage014[17]},
      {stage016[130], stage015[136], stage014[143], stage013[154], stage012[216]}
   );
   gpc615_5 gpc615_5_368(
      {stage012[113], stage012[114], stage012[115], stage012[116], stage012[117]},
      {stage013[39]},
      {stage014[18], stage014[19], stage014[20], stage014[21], stage014[22], stage014[23]},
      {stage016[131], stage015[137], stage014[144], stage013[155], stage012[217]}
   );
   gpc615_5 gpc615_5_369(
      {stage012[118], stage012[119], stage012[120], stage012[121], stage012[122]},
      {stage013[40]},
      {stage014[24], stage014[25], stage014[26], stage014[27], stage014[28], stage014[29]},
      {stage016[132], stage015[138], stage014[145], stage013[156], stage012[218]}
   );
   gpc615_5 gpc615_5_370(
      {stage012[123], stage012[124], stage012[125], stage012[126], stage012[127]},
      {stage013[41]},
      {stage014[30], stage014[31], stage014[32], stage014[33], stage014[34], stage014[35]},
      {stage016[133], stage015[139], stage014[146], stage013[157], stage012[219]}
   );
   gpc1_1 gpc1_1_371(
      {stage013[42]},
      {stage013[158]}
   );
   gpc1_1 gpc1_1_372(
      {stage013[43]},
      {stage013[159]}
   );
   gpc1_1 gpc1_1_373(
      {stage013[44]},
      {stage013[160]}
   );
   gpc1_1 gpc1_1_374(
      {stage013[45]},
      {stage013[161]}
   );
   gpc1_1 gpc1_1_375(
      {stage013[46]},
      {stage013[162]}
   );
   gpc1_1 gpc1_1_376(
      {stage013[47]},
      {stage013[163]}
   );
   gpc1_1 gpc1_1_377(
      {stage013[48]},
      {stage013[164]}
   );
   gpc1_1 gpc1_1_378(
      {stage013[49]},
      {stage013[165]}
   );
   gpc1_1 gpc1_1_379(
      {stage013[50]},
      {stage013[166]}
   );
   gpc1_1 gpc1_1_380(
      {stage013[51]},
      {stage013[167]}
   );
   gpc1_1 gpc1_1_381(
      {stage013[52]},
      {stage013[168]}
   );
   gpc1_1 gpc1_1_382(
      {stage013[53]},
      {stage013[169]}
   );
   gpc1_1 gpc1_1_383(
      {stage013[54]},
      {stage013[170]}
   );
   gpc1_1 gpc1_1_384(
      {stage013[55]},
      {stage013[171]}
   );
   gpc606_5 gpc606_5_385(
      {stage013[56], stage013[57], stage013[58], stage013[59], stage013[60], stage013[61]},
      {stage015[0], stage015[1], stage015[2], stage015[3], stage015[4], stage015[5]},
      {stage017[128], stage016[134], stage015[140], stage014[147], stage013[172]}
   );
   gpc606_5 gpc606_5_386(
      {stage013[62], stage013[63], stage013[64], stage013[65], stage013[66], stage013[67]},
      {stage015[6], stage015[7], stage015[8], stage015[9], stage015[10], stage015[11]},
      {stage017[129], stage016[135], stage015[141], stage014[148], stage013[173]}
   );
   gpc606_5 gpc606_5_387(
      {stage013[68], stage013[69], stage013[70], stage013[71], stage013[72], stage013[73]},
      {stage015[12], stage015[13], stage015[14], stage015[15], stage015[16], stage015[17]},
      {stage017[130], stage016[136], stage015[142], stage014[149], stage013[174]}
   );
   gpc606_5 gpc606_5_388(
      {stage013[74], stage013[75], stage013[76], stage013[77], stage013[78], stage013[79]},
      {stage015[18], stage015[19], stage015[20], stage015[21], stage015[22], stage015[23]},
      {stage017[131], stage016[137], stage015[143], stage014[150], stage013[175]}
   );
   gpc606_5 gpc606_5_389(
      {stage013[80], stage013[81], stage013[82], stage013[83], stage013[84], stage013[85]},
      {stage015[24], stage015[25], stage015[26], stage015[27], stage015[28], stage015[29]},
      {stage017[132], stage016[138], stage015[144], stage014[151], stage013[176]}
   );
   gpc606_5 gpc606_5_390(
      {stage013[86], stage013[87], stage013[88], stage013[89], stage013[90], stage013[91]},
      {stage015[30], stage015[31], stage015[32], stage015[33], stage015[34], stage015[35]},
      {stage017[133], stage016[139], stage015[145], stage014[152], stage013[177]}
   );
   gpc606_5 gpc606_5_391(
      {stage013[92], stage013[93], stage013[94], stage013[95], stage013[96], stage013[97]},
      {stage015[36], stage015[37], stage015[38], stage015[39], stage015[40], stage015[41]},
      {stage017[134], stage016[140], stage015[146], stage014[153], stage013[178]}
   );
   gpc606_5 gpc606_5_392(
      {stage013[98], stage013[99], stage013[100], stage013[101], stage013[102], stage013[103]},
      {stage015[42], stage015[43], stage015[44], stage015[45], stage015[46], stage015[47]},
      {stage017[135], stage016[141], stage015[147], stage014[154], stage013[179]}
   );
   gpc606_5 gpc606_5_393(
      {stage013[104], stage013[105], stage013[106], stage013[107], stage013[108], stage013[109]},
      {stage015[48], stage015[49], stage015[50], stage015[51], stage015[52], stage015[53]},
      {stage017[136], stage016[142], stage015[148], stage014[155], stage013[180]}
   );
   gpc606_5 gpc606_5_394(
      {stage013[110], stage013[111], stage013[112], stage013[113], stage013[114], stage013[115]},
      {stage015[54], stage015[55], stage015[56], stage015[57], stage015[58], stage015[59]},
      {stage017[137], stage016[143], stage015[149], stage014[156], stage013[181]}
   );
   gpc606_5 gpc606_5_395(
      {stage013[116], stage013[117], stage013[118], stage013[119], stage013[120], stage013[121]},
      {stage015[60], stage015[61], stage015[62], stage015[63], stage015[64], stage015[65]},
      {stage017[138], stage016[144], stage015[150], stage014[157], stage013[182]}
   );
   gpc606_5 gpc606_5_396(
      {stage013[122], stage013[123], stage013[124], stage013[125], stage013[126], stage013[127]},
      {stage015[66], stage015[67], stage015[68], stage015[69], stage015[70], stage015[71]},
      {stage017[139], stage016[145], stage015[151], stage014[158], stage013[183]}
   );
   gpc1_1 gpc1_1_397(
      {stage014[36]},
      {stage014[159]}
   );
   gpc1_1 gpc1_1_398(
      {stage014[37]},
      {stage014[160]}
   );
   gpc1_1 gpc1_1_399(
      {stage014[38]},
      {stage014[161]}
   );
   gpc1_1 gpc1_1_400(
      {stage014[39]},
      {stage014[162]}
   );
   gpc1_1 gpc1_1_401(
      {stage014[40]},
      {stage014[163]}
   );
   gpc1_1 gpc1_1_402(
      {stage014[41]},
      {stage014[164]}
   );
   gpc1_1 gpc1_1_403(
      {stage014[42]},
      {stage014[165]}
   );
   gpc1_1 gpc1_1_404(
      {stage014[43]},
      {stage014[166]}
   );
   gpc1_1 gpc1_1_405(
      {stage014[44]},
      {stage014[167]}
   );
   gpc1_1 gpc1_1_406(
      {stage014[45]},
      {stage014[168]}
   );
   gpc1_1 gpc1_1_407(
      {stage014[46]},
      {stage014[169]}
   );
   gpc1_1 gpc1_1_408(
      {stage014[47]},
      {stage014[170]}
   );
   gpc1_1 gpc1_1_409(
      {stage014[48]},
      {stage014[171]}
   );
   gpc1_1 gpc1_1_410(
      {stage014[49]},
      {stage014[172]}
   );
   gpc1_1 gpc1_1_411(
      {stage014[50]},
      {stage014[173]}
   );
   gpc1_1 gpc1_1_412(
      {stage014[51]},
      {stage014[174]}
   );
   gpc1_1 gpc1_1_413(
      {stage014[52]},
      {stage014[175]}
   );
   gpc1_1 gpc1_1_414(
      {stage014[53]},
      {stage014[176]}
   );
   gpc1_1 gpc1_1_415(
      {stage014[54]},
      {stage014[177]}
   );
   gpc1_1 gpc1_1_416(
      {stage014[55]},
      {stage014[178]}
   );
   gpc1_1 gpc1_1_417(
      {stage014[56]},
      {stage014[179]}
   );
   gpc1_1 gpc1_1_418(
      {stage014[57]},
      {stage014[180]}
   );
   gpc1_1 gpc1_1_419(
      {stage014[58]},
      {stage014[181]}
   );
   gpc1_1 gpc1_1_420(
      {stage014[59]},
      {stage014[182]}
   );
   gpc1_1 gpc1_1_421(
      {stage014[60]},
      {stage014[183]}
   );
   gpc1_1 gpc1_1_422(
      {stage014[61]},
      {stage014[184]}
   );
   gpc1_1 gpc1_1_423(
      {stage014[62]},
      {stage014[185]}
   );
   gpc1_1 gpc1_1_424(
      {stage014[63]},
      {stage014[186]}
   );
   gpc1_1 gpc1_1_425(
      {stage014[64]},
      {stage014[187]}
   );
   gpc1_1 gpc1_1_426(
      {stage014[65]},
      {stage014[188]}
   );
   gpc1_1 gpc1_1_427(
      {stage014[66]},
      {stage014[189]}
   );
   gpc1_1 gpc1_1_428(
      {stage014[67]},
      {stage014[190]}
   );
   gpc1_1 gpc1_1_429(
      {stage014[68]},
      {stage014[191]}
   );
   gpc1_1 gpc1_1_430(
      {stage014[69]},
      {stage014[192]}
   );
   gpc1_1 gpc1_1_431(
      {stage014[70]},
      {stage014[193]}
   );
   gpc1_1 gpc1_1_432(
      {stage014[71]},
      {stage014[194]}
   );
   gpc1_1 gpc1_1_433(
      {stage014[72]},
      {stage014[195]}
   );
   gpc1_1 gpc1_1_434(
      {stage014[73]},
      {stage014[196]}
   );
   gpc1_1 gpc1_1_435(
      {stage014[74]},
      {stage014[197]}
   );
   gpc1_1 gpc1_1_436(
      {stage014[75]},
      {stage014[198]}
   );
   gpc1_1 gpc1_1_437(
      {stage014[76]},
      {stage014[199]}
   );
   gpc1_1 gpc1_1_438(
      {stage014[77]},
      {stage014[200]}
   );
   gpc1_1 gpc1_1_439(
      {stage014[78]},
      {stage014[201]}
   );
   gpc1_1 gpc1_1_440(
      {stage014[79]},
      {stage014[202]}
   );
   gpc1_1 gpc1_1_441(
      {stage014[80]},
      {stage014[203]}
   );
   gpc1_1 gpc1_1_442(
      {stage014[81]},
      {stage014[204]}
   );
   gpc1_1 gpc1_1_443(
      {stage014[82]},
      {stage014[205]}
   );
   gpc1_1 gpc1_1_444(
      {stage014[83]},
      {stage014[206]}
   );
   gpc1_1 gpc1_1_445(
      {stage014[84]},
      {stage014[207]}
   );
   gpc1_1 gpc1_1_446(
      {stage014[85]},
      {stage014[208]}
   );
   gpc1_1 gpc1_1_447(
      {stage014[86]},
      {stage014[209]}
   );
   gpc1_1 gpc1_1_448(
      {stage014[87]},
      {stage014[210]}
   );
   gpc1_1 gpc1_1_449(
      {stage014[88]},
      {stage014[211]}
   );
   gpc1_1 gpc1_1_450(
      {stage014[89]},
      {stage014[212]}
   );
   gpc1_1 gpc1_1_451(
      {stage014[90]},
      {stage014[213]}
   );
   gpc1_1 gpc1_1_452(
      {stage014[91]},
      {stage014[214]}
   );
   gpc1_1 gpc1_1_453(
      {stage014[92]},
      {stage014[215]}
   );
   gpc1_1 gpc1_1_454(
      {stage014[93]},
      {stage014[216]}
   );
   gpc1_1 gpc1_1_455(
      {stage014[94]},
      {stage014[217]}
   );
   gpc1_1 gpc1_1_456(
      {stage014[95]},
      {stage014[218]}
   );
   gpc1_1 gpc1_1_457(
      {stage014[96]},
      {stage014[219]}
   );
   gpc1_1 gpc1_1_458(
      {stage014[97]},
      {stage014[220]}
   );
   gpc615_5 gpc615_5_459(
      {stage014[98], stage014[99], stage014[100], stage014[101], stage014[102]},
      {stage015[72]},
      {stage016[0], stage016[1], stage016[2], stage016[3], stage016[4], stage016[5]},
      {stage018[128], stage017[140], stage016[146], stage015[152], stage014[221]}
   );
   gpc615_5 gpc615_5_460(
      {stage014[103], stage014[104], stage014[105], stage014[106], stage014[107]},
      {stage015[73]},
      {stage016[6], stage016[7], stage016[8], stage016[9], stage016[10], stage016[11]},
      {stage018[129], stage017[141], stage016[147], stage015[153], stage014[222]}
   );
   gpc615_5 gpc615_5_461(
      {stage014[108], stage014[109], stage014[110], stage014[111], stage014[112]},
      {stage015[74]},
      {stage016[12], stage016[13], stage016[14], stage016[15], stage016[16], stage016[17]},
      {stage018[130], stage017[142], stage016[148], stage015[154], stage014[223]}
   );
   gpc615_5 gpc615_5_462(
      {stage014[113], stage014[114], stage014[115], stage014[116], stage014[117]},
      {stage015[75]},
      {stage016[18], stage016[19], stage016[20], stage016[21], stage016[22], stage016[23]},
      {stage018[131], stage017[143], stage016[149], stage015[155], stage014[224]}
   );
   gpc615_5 gpc615_5_463(
      {stage014[118], stage014[119], stage014[120], stage014[121], stage014[122]},
      {stage015[76]},
      {stage016[24], stage016[25], stage016[26], stage016[27], stage016[28], stage016[29]},
      {stage018[132], stage017[144], stage016[150], stage015[156], stage014[225]}
   );
   gpc615_5 gpc615_5_464(
      {stage014[123], stage014[124], stage014[125], stage014[126], stage014[127]},
      {stage015[77]},
      {stage016[30], stage016[31], stage016[32], stage016[33], stage016[34], stage016[35]},
      {stage018[133], stage017[145], stage016[151], stage015[157], stage014[226]}
   );
   gpc1_1 gpc1_1_465(
      {stage015[78]},
      {stage015[158]}
   );
   gpc1_1 gpc1_1_466(
      {stage015[79]},
      {stage015[159]}
   );
   gpc1_1 gpc1_1_467(
      {stage015[80]},
      {stage015[160]}
   );
   gpc1_1 gpc1_1_468(
      {stage015[81]},
      {stage015[161]}
   );
   gpc1_1 gpc1_1_469(
      {stage015[82]},
      {stage015[162]}
   );
   gpc1_1 gpc1_1_470(
      {stage015[83]},
      {stage015[163]}
   );
   gpc1_1 gpc1_1_471(
      {stage015[84]},
      {stage015[164]}
   );
   gpc1_1 gpc1_1_472(
      {stage015[85]},
      {stage015[165]}
   );
   gpc1_1 gpc1_1_473(
      {stage015[86]},
      {stage015[166]}
   );
   gpc1_1 gpc1_1_474(
      {stage015[87]},
      {stage015[167]}
   );
   gpc1_1 gpc1_1_475(
      {stage015[88]},
      {stage015[168]}
   );
   gpc1_1 gpc1_1_476(
      {stage015[89]},
      {stage015[169]}
   );
   gpc1_1 gpc1_1_477(
      {stage015[90]},
      {stage015[170]}
   );
   gpc1_1 gpc1_1_478(
      {stage015[91]},
      {stage015[171]}
   );
   gpc1_1 gpc1_1_479(
      {stage015[92]},
      {stage015[172]}
   );
   gpc1_1 gpc1_1_480(
      {stage015[93]},
      {stage015[173]}
   );
   gpc1_1 gpc1_1_481(
      {stage015[94]},
      {stage015[174]}
   );
   gpc1_1 gpc1_1_482(
      {stage015[95]},
      {stage015[175]}
   );
   gpc1_1 gpc1_1_483(
      {stage015[96]},
      {stage015[176]}
   );
   gpc1_1 gpc1_1_484(
      {stage015[97]},
      {stage015[177]}
   );
   gpc1_1 gpc1_1_485(
      {stage015[98]},
      {stage015[178]}
   );
   gpc1_1 gpc1_1_486(
      {stage015[99]},
      {stage015[179]}
   );
   gpc1_1 gpc1_1_487(
      {stage015[100]},
      {stage015[180]}
   );
   gpc1_1 gpc1_1_488(
      {stage015[101]},
      {stage015[181]}
   );
   gpc1_1 gpc1_1_489(
      {stage015[102]},
      {stage015[182]}
   );
   gpc615_5 gpc615_5_490(
      {stage015[103], stage015[104], stage015[105], stage015[106], stage015[107]},
      {stage016[36]},
      {stage017[0], stage017[1], stage017[2], stage017[3], stage017[4], stage017[5]},
      {stage019[128], stage018[134], stage017[146], stage016[152], stage015[183]}
   );
   gpc615_5 gpc615_5_491(
      {stage015[108], stage015[109], stage015[110], stage015[111], stage015[112]},
      {stage016[37]},
      {stage017[6], stage017[7], stage017[8], stage017[9], stage017[10], stage017[11]},
      {stage019[129], stage018[135], stage017[147], stage016[153], stage015[184]}
   );
   gpc615_5 gpc615_5_492(
      {stage015[113], stage015[114], stage015[115], stage015[116], stage015[117]},
      {stage016[38]},
      {stage017[12], stage017[13], stage017[14], stage017[15], stage017[16], stage017[17]},
      {stage019[130], stage018[136], stage017[148], stage016[154], stage015[185]}
   );
   gpc615_5 gpc615_5_493(
      {stage015[118], stage015[119], stage015[120], stage015[121], stage015[122]},
      {stage016[39]},
      {stage017[18], stage017[19], stage017[20], stage017[21], stage017[22], stage017[23]},
      {stage019[131], stage018[137], stage017[149], stage016[155], stage015[186]}
   );
   gpc615_5 gpc615_5_494(
      {stage015[123], stage015[124], stage015[125], stage015[126], stage015[127]},
      {stage016[40]},
      {stage017[24], stage017[25], stage017[26], stage017[27], stage017[28], stage017[29]},
      {stage019[132], stage018[138], stage017[150], stage016[156], stage015[187]}
   );
   gpc1_1 gpc1_1_495(
      {stage016[41]},
      {stage016[157]}
   );
   gpc1_1 gpc1_1_496(
      {stage016[42]},
      {stage016[158]}
   );
   gpc1_1 gpc1_1_497(
      {stage016[43]},
      {stage016[159]}
   );
   gpc1_1 gpc1_1_498(
      {stage016[44]},
      {stage016[160]}
   );
   gpc1_1 gpc1_1_499(
      {stage016[45]},
      {stage016[161]}
   );
   gpc1_1 gpc1_1_500(
      {stage016[46]},
      {stage016[162]}
   );
   gpc1_1 gpc1_1_501(
      {stage016[47]},
      {stage016[163]}
   );
   gpc1_1 gpc1_1_502(
      {stage016[48]},
      {stage016[164]}
   );
   gpc1_1 gpc1_1_503(
      {stage016[49]},
      {stage016[165]}
   );
   gpc1_1 gpc1_1_504(
      {stage016[50]},
      {stage016[166]}
   );
   gpc1_1 gpc1_1_505(
      {stage016[51]},
      {stage016[167]}
   );
   gpc1_1 gpc1_1_506(
      {stage016[52]},
      {stage016[168]}
   );
   gpc1_1 gpc1_1_507(
      {stage016[53]},
      {stage016[169]}
   );
   gpc1_1 gpc1_1_508(
      {stage016[54]},
      {stage016[170]}
   );
   gpc1_1 gpc1_1_509(
      {stage016[55]},
      {stage016[171]}
   );
   gpc1_1 gpc1_1_510(
      {stage016[56]},
      {stage016[172]}
   );
   gpc1_1 gpc1_1_511(
      {stage016[57]},
      {stage016[173]}
   );
   gpc1_1 gpc1_1_512(
      {stage016[58]},
      {stage016[174]}
   );
   gpc1_1 gpc1_1_513(
      {stage016[59]},
      {stage016[175]}
   );
   gpc1_1 gpc1_1_514(
      {stage016[60]},
      {stage016[176]}
   );
   gpc1_1 gpc1_1_515(
      {stage016[61]},
      {stage016[177]}
   );
   gpc1_1 gpc1_1_516(
      {stage016[62]},
      {stage016[178]}
   );
   gpc1_1 gpc1_1_517(
      {stage016[63]},
      {stage016[179]}
   );
   gpc1_1 gpc1_1_518(
      {stage016[64]},
      {stage016[180]}
   );
   gpc1_1 gpc1_1_519(
      {stage016[65]},
      {stage016[181]}
   );
   gpc1_1 gpc1_1_520(
      {stage016[66]},
      {stage016[182]}
   );
   gpc1_1 gpc1_1_521(
      {stage016[67]},
      {stage016[183]}
   );
   gpc1_1 gpc1_1_522(
      {stage016[68]},
      {stage016[184]}
   );
   gpc1_1 gpc1_1_523(
      {stage016[69]},
      {stage016[185]}
   );
   gpc1_1 gpc1_1_524(
      {stage016[70]},
      {stage016[186]}
   );
   gpc1_1 gpc1_1_525(
      {stage016[71]},
      {stage016[187]}
   );
   gpc1_1 gpc1_1_526(
      {stage016[72]},
      {stage016[188]}
   );
   gpc1_1 gpc1_1_527(
      {stage016[73]},
      {stage016[189]}
   );
   gpc1_1 gpc1_1_528(
      {stage016[74]},
      {stage016[190]}
   );
   gpc1_1 gpc1_1_529(
      {stage016[75]},
      {stage016[191]}
   );
   gpc1_1 gpc1_1_530(
      {stage016[76]},
      {stage016[192]}
   );
   gpc1_1 gpc1_1_531(
      {stage016[77]},
      {stage016[193]}
   );
   gpc1_1 gpc1_1_532(
      {stage016[78]},
      {stage016[194]}
   );
   gpc1_1 gpc1_1_533(
      {stage016[79]},
      {stage016[195]}
   );
   gpc1_1 gpc1_1_534(
      {stage016[80]},
      {stage016[196]}
   );
   gpc1_1 gpc1_1_535(
      {stage016[81]},
      {stage016[197]}
   );
   gpc1_1 gpc1_1_536(
      {stage016[82]},
      {stage016[198]}
   );
   gpc1_1 gpc1_1_537(
      {stage016[83]},
      {stage016[199]}
   );
   gpc1_1 gpc1_1_538(
      {stage016[84]},
      {stage016[200]}
   );
   gpc1_1 gpc1_1_539(
      {stage016[85]},
      {stage016[201]}
   );
   gpc606_5 gpc606_5_540(
      {stage016[86], stage016[87], stage016[88], stage016[89], stage016[90], stage016[91]},
      {stage018[0], stage018[1], stage018[2], stage018[3], stage018[4], stage018[5]},
      {stage020[128], stage019[133], stage018[139], stage017[151], stage016[202]}
   );
   gpc606_5 gpc606_5_541(
      {stage016[92], stage016[93], stage016[94], stage016[95], stage016[96], stage016[97]},
      {stage018[6], stage018[7], stage018[8], stage018[9], stage018[10], stage018[11]},
      {stage020[129], stage019[134], stage018[140], stage017[152], stage016[203]}
   );
   gpc606_5 gpc606_5_542(
      {stage016[98], stage016[99], stage016[100], stage016[101], stage016[102], stage016[103]},
      {stage018[12], stage018[13], stage018[14], stage018[15], stage018[16], stage018[17]},
      {stage020[130], stage019[135], stage018[141], stage017[153], stage016[204]}
   );
   gpc606_5 gpc606_5_543(
      {stage016[104], stage016[105], stage016[106], stage016[107], stage016[108], stage016[109]},
      {stage018[18], stage018[19], stage018[20], stage018[21], stage018[22], stage018[23]},
      {stage020[131], stage019[136], stage018[142], stage017[154], stage016[205]}
   );
   gpc606_5 gpc606_5_544(
      {stage016[110], stage016[111], stage016[112], stage016[113], stage016[114], stage016[115]},
      {stage018[24], stage018[25], stage018[26], stage018[27], stage018[28], stage018[29]},
      {stage020[132], stage019[137], stage018[143], stage017[155], stage016[206]}
   );
   gpc606_5 gpc606_5_545(
      {stage016[116], stage016[117], stage016[118], stage016[119], stage016[120], stage016[121]},
      {stage018[30], stage018[31], stage018[32], stage018[33], stage018[34], stage018[35]},
      {stage020[133], stage019[138], stage018[144], stage017[156], stage016[207]}
   );
   gpc606_5 gpc606_5_546(
      {stage016[122], stage016[123], stage016[124], stage016[125], stage016[126], stage016[127]},
      {stage018[36], stage018[37], stage018[38], stage018[39], stage018[40], stage018[41]},
      {stage020[134], stage019[139], stage018[145], stage017[157], stage016[208]}
   );
   gpc1_1 gpc1_1_547(
      {stage017[30]},
      {stage017[158]}
   );
   gpc1_1 gpc1_1_548(
      {stage017[31]},
      {stage017[159]}
   );
   gpc1_1 gpc1_1_549(
      {stage017[32]},
      {stage017[160]}
   );
   gpc1_1 gpc1_1_550(
      {stage017[33]},
      {stage017[161]}
   );
   gpc1_1 gpc1_1_551(
      {stage017[34]},
      {stage017[162]}
   );
   gpc1_1 gpc1_1_552(
      {stage017[35]},
      {stage017[163]}
   );
   gpc1_1 gpc1_1_553(
      {stage017[36]},
      {stage017[164]}
   );
   gpc1_1 gpc1_1_554(
      {stage017[37]},
      {stage017[165]}
   );
   gpc1_1 gpc1_1_555(
      {stage017[38]},
      {stage017[166]}
   );
   gpc1_1 gpc1_1_556(
      {stage017[39]},
      {stage017[167]}
   );
   gpc1_1 gpc1_1_557(
      {stage017[40]},
      {stage017[168]}
   );
   gpc1_1 gpc1_1_558(
      {stage017[41]},
      {stage017[169]}
   );
   gpc1_1 gpc1_1_559(
      {stage017[42]},
      {stage017[170]}
   );
   gpc1_1 gpc1_1_560(
      {stage017[43]},
      {stage017[171]}
   );
   gpc1_1 gpc1_1_561(
      {stage017[44]},
      {stage017[172]}
   );
   gpc1_1 gpc1_1_562(
      {stage017[45]},
      {stage017[173]}
   );
   gpc1_1 gpc1_1_563(
      {stage017[46]},
      {stage017[174]}
   );
   gpc1_1 gpc1_1_564(
      {stage017[47]},
      {stage017[175]}
   );
   gpc1_1 gpc1_1_565(
      {stage017[48]},
      {stage017[176]}
   );
   gpc1_1 gpc1_1_566(
      {stage017[49]},
      {stage017[177]}
   );
   gpc1_1 gpc1_1_567(
      {stage017[50]},
      {stage017[178]}
   );
   gpc1_1 gpc1_1_568(
      {stage017[51]},
      {stage017[179]}
   );
   gpc1_1 gpc1_1_569(
      {stage017[52]},
      {stage017[180]}
   );
   gpc1_1 gpc1_1_570(
      {stage017[53]},
      {stage017[181]}
   );
   gpc1_1 gpc1_1_571(
      {stage017[54]},
      {stage017[182]}
   );
   gpc1_1 gpc1_1_572(
      {stage017[55]},
      {stage017[183]}
   );
   gpc1_1 gpc1_1_573(
      {stage017[56]},
      {stage017[184]}
   );
   gpc1_1 gpc1_1_574(
      {stage017[57]},
      {stage017[185]}
   );
   gpc1_1 gpc1_1_575(
      {stage017[58]},
      {stage017[186]}
   );
   gpc1_1 gpc1_1_576(
      {stage017[59]},
      {stage017[187]}
   );
   gpc1_1 gpc1_1_577(
      {stage017[60]},
      {stage017[188]}
   );
   gpc1_1 gpc1_1_578(
      {stage017[61]},
      {stage017[189]}
   );
   gpc1_1 gpc1_1_579(
      {stage017[62]},
      {stage017[190]}
   );
   gpc1_1 gpc1_1_580(
      {stage017[63]},
      {stage017[191]}
   );
   gpc1_1 gpc1_1_581(
      {stage017[64]},
      {stage017[192]}
   );
   gpc1_1 gpc1_1_582(
      {stage017[65]},
      {stage017[193]}
   );
   gpc1_1 gpc1_1_583(
      {stage017[66]},
      {stage017[194]}
   );
   gpc1_1 gpc1_1_584(
      {stage017[67]},
      {stage017[195]}
   );
   gpc1_1 gpc1_1_585(
      {stage017[68]},
      {stage017[196]}
   );
   gpc1_1 gpc1_1_586(
      {stage017[69]},
      {stage017[197]}
   );
   gpc1_1 gpc1_1_587(
      {stage017[70]},
      {stage017[198]}
   );
   gpc1_1 gpc1_1_588(
      {stage017[71]},
      {stage017[199]}
   );
   gpc1_1 gpc1_1_589(
      {stage017[72]},
      {stage017[200]}
   );
   gpc1_1 gpc1_1_590(
      {stage017[73]},
      {stage017[201]}
   );
   gpc1_1 gpc1_1_591(
      {stage017[74]},
      {stage017[202]}
   );
   gpc1_1 gpc1_1_592(
      {stage017[75]},
      {stage017[203]}
   );
   gpc1_1 gpc1_1_593(
      {stage017[76]},
      {stage017[204]}
   );
   gpc1_1 gpc1_1_594(
      {stage017[77]},
      {stage017[205]}
   );
   gpc1_1 gpc1_1_595(
      {stage017[78]},
      {stage017[206]}
   );
   gpc1_1 gpc1_1_596(
      {stage017[79]},
      {stage017[207]}
   );
   gpc1_1 gpc1_1_597(
      {stage017[80]},
      {stage017[208]}
   );
   gpc1_1 gpc1_1_598(
      {stage017[81]},
      {stage017[209]}
   );
   gpc606_5 gpc606_5_599(
      {stage017[82], stage017[83], stage017[84], stage017[85], stage017[86], stage017[87]},
      {stage019[0], stage019[1], stage019[2], stage019[3], stage019[4], stage019[5]},
      {stage021[128], stage020[135], stage019[140], stage018[146], stage017[210]}
   );
   gpc615_5 gpc615_5_600(
      {stage017[88], stage017[89], stage017[90], stage017[91], stage017[92]},
      {stage018[42]},
      {stage019[6], stage019[7], stage019[8], stage019[9], stage019[10], stage019[11]},
      {stage021[129], stage020[136], stage019[141], stage018[147], stage017[211]}
   );
   gpc615_5 gpc615_5_601(
      {stage017[93], stage017[94], stage017[95], stage017[96], stage017[97]},
      {stage018[43]},
      {stage019[12], stage019[13], stage019[14], stage019[15], stage019[16], stage019[17]},
      {stage021[130], stage020[137], stage019[142], stage018[148], stage017[212]}
   );
   gpc615_5 gpc615_5_602(
      {stage017[98], stage017[99], stage017[100], stage017[101], stage017[102]},
      {stage018[44]},
      {stage019[18], stage019[19], stage019[20], stage019[21], stage019[22], stage019[23]},
      {stage021[131], stage020[138], stage019[143], stage018[149], stage017[213]}
   );
   gpc615_5 gpc615_5_603(
      {stage017[103], stage017[104], stage017[105], stage017[106], stage017[107]},
      {stage018[45]},
      {stage019[24], stage019[25], stage019[26], stage019[27], stage019[28], stage019[29]},
      {stage021[132], stage020[139], stage019[144], stage018[150], stage017[214]}
   );
   gpc615_5 gpc615_5_604(
      {stage017[108], stage017[109], stage017[110], stage017[111], stage017[112]},
      {stage018[46]},
      {stage019[30], stage019[31], stage019[32], stage019[33], stage019[34], stage019[35]},
      {stage021[133], stage020[140], stage019[145], stage018[151], stage017[215]}
   );
   gpc615_5 gpc615_5_605(
      {stage017[113], stage017[114], stage017[115], stage017[116], stage017[117]},
      {stage018[47]},
      {stage019[36], stage019[37], stage019[38], stage019[39], stage019[40], stage019[41]},
      {stage021[134], stage020[141], stage019[146], stage018[152], stage017[216]}
   );
   gpc615_5 gpc615_5_606(
      {stage017[118], stage017[119], stage017[120], stage017[121], stage017[122]},
      {stage018[48]},
      {stage019[42], stage019[43], stage019[44], stage019[45], stage019[46], stage019[47]},
      {stage021[135], stage020[142], stage019[147], stage018[153], stage017[217]}
   );
   gpc615_5 gpc615_5_607(
      {stage017[123], stage017[124], stage017[125], stage017[126], stage017[127]},
      {stage018[49]},
      {stage019[48], stage019[49], stage019[50], stage019[51], stage019[52], stage019[53]},
      {stage021[136], stage020[143], stage019[148], stage018[154], stage017[218]}
   );
   gpc1_1 gpc1_1_608(
      {stage018[50]},
      {stage018[155]}
   );
   gpc1_1 gpc1_1_609(
      {stage018[51]},
      {stage018[156]}
   );
   gpc1_1 gpc1_1_610(
      {stage018[52]},
      {stage018[157]}
   );
   gpc1_1 gpc1_1_611(
      {stage018[53]},
      {stage018[158]}
   );
   gpc1_1 gpc1_1_612(
      {stage018[54]},
      {stage018[159]}
   );
   gpc1_1 gpc1_1_613(
      {stage018[55]},
      {stage018[160]}
   );
   gpc1_1 gpc1_1_614(
      {stage018[56]},
      {stage018[161]}
   );
   gpc1_1 gpc1_1_615(
      {stage018[57]},
      {stage018[162]}
   );
   gpc1_1 gpc1_1_616(
      {stage018[58]},
      {stage018[163]}
   );
   gpc1_1 gpc1_1_617(
      {stage018[59]},
      {stage018[164]}
   );
   gpc1_1 gpc1_1_618(
      {stage018[60]},
      {stage018[165]}
   );
   gpc1_1 gpc1_1_619(
      {stage018[61]},
      {stage018[166]}
   );
   gpc1_1 gpc1_1_620(
      {stage018[62]},
      {stage018[167]}
   );
   gpc1_1 gpc1_1_621(
      {stage018[63]},
      {stage018[168]}
   );
   gpc1_1 gpc1_1_622(
      {stage018[64]},
      {stage018[169]}
   );
   gpc1_1 gpc1_1_623(
      {stage018[65]},
      {stage018[170]}
   );
   gpc1_1 gpc1_1_624(
      {stage018[66]},
      {stage018[171]}
   );
   gpc1_1 gpc1_1_625(
      {stage018[67]},
      {stage018[172]}
   );
   gpc1_1 gpc1_1_626(
      {stage018[68]},
      {stage018[173]}
   );
   gpc1_1 gpc1_1_627(
      {stage018[69]},
      {stage018[174]}
   );
   gpc1_1 gpc1_1_628(
      {stage018[70]},
      {stage018[175]}
   );
   gpc1_1 gpc1_1_629(
      {stage018[71]},
      {stage018[176]}
   );
   gpc1_1 gpc1_1_630(
      {stage018[72]},
      {stage018[177]}
   );
   gpc615_5 gpc615_5_631(
      {stage018[73], stage018[74], stage018[75], stage018[76], stage018[77]},
      {stage019[54]},
      {stage020[0], stage020[1], stage020[2], stage020[3], stage020[4], stage020[5]},
      {stage022[128], stage021[137], stage020[144], stage019[149], stage018[178]}
   );
   gpc615_5 gpc615_5_632(
      {stage018[78], stage018[79], stage018[80], stage018[81], stage018[82]},
      {stage019[55]},
      {stage020[6], stage020[7], stage020[8], stage020[9], stage020[10], stage020[11]},
      {stage022[129], stage021[138], stage020[145], stage019[150], stage018[179]}
   );
   gpc615_5 gpc615_5_633(
      {stage018[83], stage018[84], stage018[85], stage018[86], stage018[87]},
      {stage019[56]},
      {stage020[12], stage020[13], stage020[14], stage020[15], stage020[16], stage020[17]},
      {stage022[130], stage021[139], stage020[146], stage019[151], stage018[180]}
   );
   gpc615_5 gpc615_5_634(
      {stage018[88], stage018[89], stage018[90], stage018[91], stage018[92]},
      {stage019[57]},
      {stage020[18], stage020[19], stage020[20], stage020[21], stage020[22], stage020[23]},
      {stage022[131], stage021[140], stage020[147], stage019[152], stage018[181]}
   );
   gpc615_5 gpc615_5_635(
      {stage018[93], stage018[94], stage018[95], stage018[96], stage018[97]},
      {stage019[58]},
      {stage020[24], stage020[25], stage020[26], stage020[27], stage020[28], stage020[29]},
      {stage022[132], stage021[141], stage020[148], stage019[153], stage018[182]}
   );
   gpc615_5 gpc615_5_636(
      {stage018[98], stage018[99], stage018[100], stage018[101], stage018[102]},
      {stage019[59]},
      {stage020[30], stage020[31], stage020[32], stage020[33], stage020[34], stage020[35]},
      {stage022[133], stage021[142], stage020[149], stage019[154], stage018[183]}
   );
   gpc615_5 gpc615_5_637(
      {stage018[103], stage018[104], stage018[105], stage018[106], stage018[107]},
      {stage019[60]},
      {stage020[36], stage020[37], stage020[38], stage020[39], stage020[40], stage020[41]},
      {stage022[134], stage021[143], stage020[150], stage019[155], stage018[184]}
   );
   gpc615_5 gpc615_5_638(
      {stage018[108], stage018[109], stage018[110], stage018[111], stage018[112]},
      {stage019[61]},
      {stage020[42], stage020[43], stage020[44], stage020[45], stage020[46], stage020[47]},
      {stage022[135], stage021[144], stage020[151], stage019[156], stage018[185]}
   );
   gpc615_5 gpc615_5_639(
      {stage018[113], stage018[114], stage018[115], stage018[116], stage018[117]},
      {stage019[62]},
      {stage020[48], stage020[49], stage020[50], stage020[51], stage020[52], stage020[53]},
      {stage022[136], stage021[145], stage020[152], stage019[157], stage018[186]}
   );
   gpc615_5 gpc615_5_640(
      {stage018[118], stage018[119], stage018[120], stage018[121], stage018[122]},
      {stage019[63]},
      {stage020[54], stage020[55], stage020[56], stage020[57], stage020[58], stage020[59]},
      {stage022[137], stage021[146], stage020[153], stage019[158], stage018[187]}
   );
   gpc615_5 gpc615_5_641(
      {stage018[123], stage018[124], stage018[125], stage018[126], stage018[127]},
      {stage019[64]},
      {stage020[60], stage020[61], stage020[62], stage020[63], stage020[64], stage020[65]},
      {stage022[138], stage021[147], stage020[154], stage019[159], stage018[188]}
   );
   gpc1_1 gpc1_1_642(
      {stage019[65]},
      {stage019[160]}
   );
   gpc1_1 gpc1_1_643(
      {stage019[66]},
      {stage019[161]}
   );
   gpc1_1 gpc1_1_644(
      {stage019[67]},
      {stage019[162]}
   );
   gpc1_1 gpc1_1_645(
      {stage019[68]},
      {stage019[163]}
   );
   gpc1_1 gpc1_1_646(
      {stage019[69]},
      {stage019[164]}
   );
   gpc1_1 gpc1_1_647(
      {stage019[70]},
      {stage019[165]}
   );
   gpc1_1 gpc1_1_648(
      {stage019[71]},
      {stage019[166]}
   );
   gpc1_1 gpc1_1_649(
      {stage019[72]},
      {stage019[167]}
   );
   gpc1_1 gpc1_1_650(
      {stage019[73]},
      {stage019[168]}
   );
   gpc1_1 gpc1_1_651(
      {stage019[74]},
      {stage019[169]}
   );
   gpc1_1 gpc1_1_652(
      {stage019[75]},
      {stage019[170]}
   );
   gpc1_1 gpc1_1_653(
      {stage019[76]},
      {stage019[171]}
   );
   gpc1_1 gpc1_1_654(
      {stage019[77]},
      {stage019[172]}
   );
   gpc1_1 gpc1_1_655(
      {stage019[78]},
      {stage019[173]}
   );
   gpc1_1 gpc1_1_656(
      {stage019[79]},
      {stage019[174]}
   );
   gpc1_1 gpc1_1_657(
      {stage019[80]},
      {stage019[175]}
   );
   gpc1_1 gpc1_1_658(
      {stage019[81]},
      {stage019[176]}
   );
   gpc1_1 gpc1_1_659(
      {stage019[82]},
      {stage019[177]}
   );
   gpc1_1 gpc1_1_660(
      {stage019[83]},
      {stage019[178]}
   );
   gpc1_1 gpc1_1_661(
      {stage019[84]},
      {stage019[179]}
   );
   gpc1_1 gpc1_1_662(
      {stage019[85]},
      {stage019[180]}
   );
   gpc606_5 gpc606_5_663(
      {stage019[86], stage019[87], stage019[88], stage019[89], stage019[90], stage019[91]},
      {stage021[0], stage021[1], stage021[2], stage021[3], stage021[4], stage021[5]},
      {stage023[128], stage022[139], stage021[148], stage020[155], stage019[181]}
   );
   gpc606_5 gpc606_5_664(
      {stage019[92], stage019[93], stage019[94], stage019[95], stage019[96], stage019[97]},
      {stage021[6], stage021[7], stage021[8], stage021[9], stage021[10], stage021[11]},
      {stage023[129], stage022[140], stage021[149], stage020[156], stage019[182]}
   );
   gpc606_5 gpc606_5_665(
      {stage019[98], stage019[99], stage019[100], stage019[101], stage019[102], stage019[103]},
      {stage021[12], stage021[13], stage021[14], stage021[15], stage021[16], stage021[17]},
      {stage023[130], stage022[141], stage021[150], stage020[157], stage019[183]}
   );
   gpc606_5 gpc606_5_666(
      {stage019[104], stage019[105], stage019[106], stage019[107], stage019[108], stage019[109]},
      {stage021[18], stage021[19], stage021[20], stage021[21], stage021[22], stage021[23]},
      {stage023[131], stage022[142], stage021[151], stage020[158], stage019[184]}
   );
   gpc606_5 gpc606_5_667(
      {stage019[110], stage019[111], stage019[112], stage019[113], stage019[114], stage019[115]},
      {stage021[24], stage021[25], stage021[26], stage021[27], stage021[28], stage021[29]},
      {stage023[132], stage022[143], stage021[152], stage020[159], stage019[185]}
   );
   gpc606_5 gpc606_5_668(
      {stage019[116], stage019[117], stage019[118], stage019[119], stage019[120], stage019[121]},
      {stage021[30], stage021[31], stage021[32], stage021[33], stage021[34], stage021[35]},
      {stage023[133], stage022[144], stage021[153], stage020[160], stage019[186]}
   );
   gpc606_5 gpc606_5_669(
      {stage019[122], stage019[123], stage019[124], stage019[125], stage019[126], stage019[127]},
      {stage021[36], stage021[37], stage021[38], stage021[39], stage021[40], stage021[41]},
      {stage023[134], stage022[145], stage021[154], stage020[161], stage019[187]}
   );
   gpc1_1 gpc1_1_670(
      {stage020[66]},
      {stage020[162]}
   );
   gpc1_1 gpc1_1_671(
      {stage020[67]},
      {stage020[163]}
   );
   gpc1_1 gpc1_1_672(
      {stage020[68]},
      {stage020[164]}
   );
   gpc1_1 gpc1_1_673(
      {stage020[69]},
      {stage020[165]}
   );
   gpc1_1 gpc1_1_674(
      {stage020[70]},
      {stage020[166]}
   );
   gpc1_1 gpc1_1_675(
      {stage020[71]},
      {stage020[167]}
   );
   gpc1_1 gpc1_1_676(
      {stage020[72]},
      {stage020[168]}
   );
   gpc1_1 gpc1_1_677(
      {stage020[73]},
      {stage020[169]}
   );
   gpc1_1 gpc1_1_678(
      {stage020[74]},
      {stage020[170]}
   );
   gpc1_1 gpc1_1_679(
      {stage020[75]},
      {stage020[171]}
   );
   gpc1_1 gpc1_1_680(
      {stage020[76]},
      {stage020[172]}
   );
   gpc1_1 gpc1_1_681(
      {stage020[77]},
      {stage020[173]}
   );
   gpc615_5 gpc615_5_682(
      {stage020[78], stage020[79], stage020[80], stage020[81], stage020[82]},
      {stage021[42]},
      {stage022[0], stage022[1], stage022[2], stage022[3], stage022[4], stage022[5]},
      {stage024[128], stage023[135], stage022[146], stage021[155], stage020[174]}
   );
   gpc615_5 gpc615_5_683(
      {stage020[83], stage020[84], stage020[85], stage020[86], stage020[87]},
      {stage021[43]},
      {stage022[6], stage022[7], stage022[8], stage022[9], stage022[10], stage022[11]},
      {stage024[129], stage023[136], stage022[147], stage021[156], stage020[175]}
   );
   gpc615_5 gpc615_5_684(
      {stage020[88], stage020[89], stage020[90], stage020[91], stage020[92]},
      {stage021[44]},
      {stage022[12], stage022[13], stage022[14], stage022[15], stage022[16], stage022[17]},
      {stage024[130], stage023[137], stage022[148], stage021[157], stage020[176]}
   );
   gpc615_5 gpc615_5_685(
      {stage020[93], stage020[94], stage020[95], stage020[96], stage020[97]},
      {stage021[45]},
      {stage022[18], stage022[19], stage022[20], stage022[21], stage022[22], stage022[23]},
      {stage024[131], stage023[138], stage022[149], stage021[158], stage020[177]}
   );
   gpc615_5 gpc615_5_686(
      {stage020[98], stage020[99], stage020[100], stage020[101], stage020[102]},
      {stage021[46]},
      {stage022[24], stage022[25], stage022[26], stage022[27], stage022[28], stage022[29]},
      {stage024[132], stage023[139], stage022[150], stage021[159], stage020[178]}
   );
   gpc615_5 gpc615_5_687(
      {stage020[103], stage020[104], stage020[105], stage020[106], stage020[107]},
      {stage021[47]},
      {stage022[30], stage022[31], stage022[32], stage022[33], stage022[34], stage022[35]},
      {stage024[133], stage023[140], stage022[151], stage021[160], stage020[179]}
   );
   gpc615_5 gpc615_5_688(
      {stage020[108], stage020[109], stage020[110], stage020[111], stage020[112]},
      {stage021[48]},
      {stage022[36], stage022[37], stage022[38], stage022[39], stage022[40], stage022[41]},
      {stage024[134], stage023[141], stage022[152], stage021[161], stage020[180]}
   );
   gpc615_5 gpc615_5_689(
      {stage020[113], stage020[114], stage020[115], stage020[116], stage020[117]},
      {stage021[49]},
      {stage022[42], stage022[43], stage022[44], stage022[45], stage022[46], stage022[47]},
      {stage024[135], stage023[142], stage022[153], stage021[162], stage020[181]}
   );
   gpc615_5 gpc615_5_690(
      {stage020[118], stage020[119], stage020[120], stage020[121], stage020[122]},
      {stage021[50]},
      {stage022[48], stage022[49], stage022[50], stage022[51], stage022[52], stage022[53]},
      {stage024[136], stage023[143], stage022[154], stage021[163], stage020[182]}
   );
   gpc615_5 gpc615_5_691(
      {stage020[123], stage020[124], stage020[125], stage020[126], stage020[127]},
      {stage021[51]},
      {stage022[54], stage022[55], stage022[56], stage022[57], stage022[58], stage022[59]},
      {stage024[137], stage023[144], stage022[155], stage021[164], stage020[183]}
   );
   gpc1_1 gpc1_1_692(
      {stage021[52]},
      {stage021[165]}
   );
   gpc1_1 gpc1_1_693(
      {stage021[53]},
      {stage021[166]}
   );
   gpc1_1 gpc1_1_694(
      {stage021[54]},
      {stage021[167]}
   );
   gpc1_1 gpc1_1_695(
      {stage021[55]},
      {stage021[168]}
   );
   gpc1_1 gpc1_1_696(
      {stage021[56]},
      {stage021[169]}
   );
   gpc1_1 gpc1_1_697(
      {stage021[57]},
      {stage021[170]}
   );
   gpc1_1 gpc1_1_698(
      {stage021[58]},
      {stage021[171]}
   );
   gpc1_1 gpc1_1_699(
      {stage021[59]},
      {stage021[172]}
   );
   gpc1_1 gpc1_1_700(
      {stage021[60]},
      {stage021[173]}
   );
   gpc1_1 gpc1_1_701(
      {stage021[61]},
      {stage021[174]}
   );
   gpc1_1 gpc1_1_702(
      {stage021[62]},
      {stage021[175]}
   );
   gpc1_1 gpc1_1_703(
      {stage021[63]},
      {stage021[176]}
   );
   gpc1_1 gpc1_1_704(
      {stage021[64]},
      {stage021[177]}
   );
   gpc1_1 gpc1_1_705(
      {stage021[65]},
      {stage021[178]}
   );
   gpc1_1 gpc1_1_706(
      {stage021[66]},
      {stage021[179]}
   );
   gpc1_1 gpc1_1_707(
      {stage021[67]},
      {stage021[180]}
   );
   gpc1_1 gpc1_1_708(
      {stage021[68]},
      {stage021[181]}
   );
   gpc1_1 gpc1_1_709(
      {stage021[69]},
      {stage021[182]}
   );
   gpc1_1 gpc1_1_710(
      {stage021[70]},
      {stage021[183]}
   );
   gpc1_1 gpc1_1_711(
      {stage021[71]},
      {stage021[184]}
   );
   gpc1_1 gpc1_1_712(
      {stage021[72]},
      {stage021[185]}
   );
   gpc1_1 gpc1_1_713(
      {stage021[73]},
      {stage021[186]}
   );
   gpc1_1 gpc1_1_714(
      {stage021[74]},
      {stage021[187]}
   );
   gpc1_1 gpc1_1_715(
      {stage021[75]},
      {stage021[188]}
   );
   gpc1_1 gpc1_1_716(
      {stage021[76]},
      {stage021[189]}
   );
   gpc1_1 gpc1_1_717(
      {stage021[77]},
      {stage021[190]}
   );
   gpc615_5 gpc615_5_718(
      {stage021[78], stage021[79], stage021[80], stage021[81], stage021[82]},
      {stage022[60]},
      {stage023[0], stage023[1], stage023[2], stage023[3], stage023[4], stage023[5]},
      {stage025[128], stage024[138], stage023[145], stage022[156], stage021[191]}
   );
   gpc615_5 gpc615_5_719(
      {stage021[83], stage021[84], stage021[85], stage021[86], stage021[87]},
      {stage022[61]},
      {stage023[6], stage023[7], stage023[8], stage023[9], stage023[10], stage023[11]},
      {stage025[129], stage024[139], stage023[146], stage022[157], stage021[192]}
   );
   gpc615_5 gpc615_5_720(
      {stage021[88], stage021[89], stage021[90], stage021[91], stage021[92]},
      {stage022[62]},
      {stage023[12], stage023[13], stage023[14], stage023[15], stage023[16], stage023[17]},
      {stage025[130], stage024[140], stage023[147], stage022[158], stage021[193]}
   );
   gpc615_5 gpc615_5_721(
      {stage021[93], stage021[94], stage021[95], stage021[96], stage021[97]},
      {stage022[63]},
      {stage023[18], stage023[19], stage023[20], stage023[21], stage023[22], stage023[23]},
      {stage025[131], stage024[141], stage023[148], stage022[159], stage021[194]}
   );
   gpc615_5 gpc615_5_722(
      {stage021[98], stage021[99], stage021[100], stage021[101], stage021[102]},
      {stage022[64]},
      {stage023[24], stage023[25], stage023[26], stage023[27], stage023[28], stage023[29]},
      {stage025[132], stage024[142], stage023[149], stage022[160], stage021[195]}
   );
   gpc615_5 gpc615_5_723(
      {stage021[103], stage021[104], stage021[105], stage021[106], stage021[107]},
      {stage022[65]},
      {stage023[30], stage023[31], stage023[32], stage023[33], stage023[34], stage023[35]},
      {stage025[133], stage024[143], stage023[150], stage022[161], stage021[196]}
   );
   gpc615_5 gpc615_5_724(
      {stage021[108], stage021[109], stage021[110], stage021[111], stage021[112]},
      {stage022[66]},
      {stage023[36], stage023[37], stage023[38], stage023[39], stage023[40], stage023[41]},
      {stage025[134], stage024[144], stage023[151], stage022[162], stage021[197]}
   );
   gpc615_5 gpc615_5_725(
      {stage021[113], stage021[114], stage021[115], stage021[116], stage021[117]},
      {stage022[67]},
      {stage023[42], stage023[43], stage023[44], stage023[45], stage023[46], stage023[47]},
      {stage025[135], stage024[145], stage023[152], stage022[163], stage021[198]}
   );
   gpc615_5 gpc615_5_726(
      {stage021[118], stage021[119], stage021[120], stage021[121], stage021[122]},
      {stage022[68]},
      {stage023[48], stage023[49], stage023[50], stage023[51], stage023[52], stage023[53]},
      {stage025[136], stage024[146], stage023[153], stage022[164], stage021[199]}
   );
   gpc615_5 gpc615_5_727(
      {stage021[123], stage021[124], stage021[125], stage021[126], stage021[127]},
      {stage022[69]},
      {stage023[54], stage023[55], stage023[56], stage023[57], stage023[58], stage023[59]},
      {stage025[137], stage024[147], stage023[154], stage022[165], stage021[200]}
   );
   gpc1_1 gpc1_1_728(
      {stage022[70]},
      {stage022[166]}
   );
   gpc1_1 gpc1_1_729(
      {stage022[71]},
      {stage022[167]}
   );
   gpc1_1 gpc1_1_730(
      {stage022[72]},
      {stage022[168]}
   );
   gpc1_1 gpc1_1_731(
      {stage022[73]},
      {stage022[169]}
   );
   gpc606_5 gpc606_5_732(
      {stage022[74], stage022[75], stage022[76], stage022[77], stage022[78], stage022[79]},
      {stage024[0], stage024[1], stage024[2], stage024[3], stage024[4], stage024[5]},
      {stage026[128], stage025[138], stage024[148], stage023[155], stage022[170]}
   );
   gpc606_5 gpc606_5_733(
      {stage022[80], stage022[81], stage022[82], stage022[83], stage022[84], stage022[85]},
      {stage024[6], stage024[7], stage024[8], stage024[9], stage024[10], stage024[11]},
      {stage026[129], stage025[139], stage024[149], stage023[156], stage022[171]}
   );
   gpc606_5 gpc606_5_734(
      {stage022[86], stage022[87], stage022[88], stage022[89], stage022[90], stage022[91]},
      {stage024[12], stage024[13], stage024[14], stage024[15], stage024[16], stage024[17]},
      {stage026[130], stage025[140], stage024[150], stage023[157], stage022[172]}
   );
   gpc606_5 gpc606_5_735(
      {stage022[92], stage022[93], stage022[94], stage022[95], stage022[96], stage022[97]},
      {stage024[18], stage024[19], stage024[20], stage024[21], stage024[22], stage024[23]},
      {stage026[131], stage025[141], stage024[151], stage023[158], stage022[173]}
   );
   gpc615_5 gpc615_5_736(
      {stage022[98], stage022[99], stage022[100], stage022[101], stage022[102]},
      {stage023[60]},
      {stage024[24], stage024[25], stage024[26], stage024[27], stage024[28], stage024[29]},
      {stage026[132], stage025[142], stage024[152], stage023[159], stage022[174]}
   );
   gpc615_5 gpc615_5_737(
      {stage022[103], stage022[104], stage022[105], stage022[106], stage022[107]},
      {stage023[61]},
      {stage024[30], stage024[31], stage024[32], stage024[33], stage024[34], stage024[35]},
      {stage026[133], stage025[143], stage024[153], stage023[160], stage022[175]}
   );
   gpc615_5 gpc615_5_738(
      {stage022[108], stage022[109], stage022[110], stage022[111], stage022[112]},
      {stage023[62]},
      {stage024[36], stage024[37], stage024[38], stage024[39], stage024[40], stage024[41]},
      {stage026[134], stage025[144], stage024[154], stage023[161], stage022[176]}
   );
   gpc615_5 gpc615_5_739(
      {stage022[113], stage022[114], stage022[115], stage022[116], stage022[117]},
      {stage023[63]},
      {stage024[42], stage024[43], stage024[44], stage024[45], stage024[46], stage024[47]},
      {stage026[135], stage025[145], stage024[155], stage023[162], stage022[177]}
   );
   gpc615_5 gpc615_5_740(
      {stage022[118], stage022[119], stage022[120], stage022[121], stage022[122]},
      {stage023[64]},
      {stage024[48], stage024[49], stage024[50], stage024[51], stage024[52], stage024[53]},
      {stage026[136], stage025[146], stage024[156], stage023[163], stage022[178]}
   );
   gpc615_5 gpc615_5_741(
      {stage022[123], stage022[124], stage022[125], stage022[126], stage022[127]},
      {stage023[65]},
      {stage024[54], stage024[55], stage024[56], stage024[57], stage024[58], stage024[59]},
      {stage026[137], stage025[147], stage024[157], stage023[164], stage022[179]}
   );
   gpc1_1 gpc1_1_742(
      {stage023[66]},
      {stage023[165]}
   );
   gpc1_1 gpc1_1_743(
      {stage023[67]},
      {stage023[166]}
   );
   gpc1_1 gpc1_1_744(
      {stage023[68]},
      {stage023[167]}
   );
   gpc1_1 gpc1_1_745(
      {stage023[69]},
      {stage023[168]}
   );
   gpc1_1 gpc1_1_746(
      {stage023[70]},
      {stage023[169]}
   );
   gpc1_1 gpc1_1_747(
      {stage023[71]},
      {stage023[170]}
   );
   gpc1_1 gpc1_1_748(
      {stage023[72]},
      {stage023[171]}
   );
   gpc1_1 gpc1_1_749(
      {stage023[73]},
      {stage023[172]}
   );
   gpc1_1 gpc1_1_750(
      {stage023[74]},
      {stage023[173]}
   );
   gpc1_1 gpc1_1_751(
      {stage023[75]},
      {stage023[174]}
   );
   gpc1_1 gpc1_1_752(
      {stage023[76]},
      {stage023[175]}
   );
   gpc1_1 gpc1_1_753(
      {stage023[77]},
      {stage023[176]}
   );
   gpc1_1 gpc1_1_754(
      {stage023[78]},
      {stage023[177]}
   );
   gpc1_1 gpc1_1_755(
      {stage023[79]},
      {stage023[178]}
   );
   gpc1_1 gpc1_1_756(
      {stage023[80]},
      {stage023[179]}
   );
   gpc1_1 gpc1_1_757(
      {stage023[81]},
      {stage023[180]}
   );
   gpc1_1 gpc1_1_758(
      {stage023[82]},
      {stage023[181]}
   );
   gpc1_1 gpc1_1_759(
      {stage023[83]},
      {stage023[182]}
   );
   gpc1_1 gpc1_1_760(
      {stage023[84]},
      {stage023[183]}
   );
   gpc1_1 gpc1_1_761(
      {stage023[85]},
      {stage023[184]}
   );
   gpc1_1 gpc1_1_762(
      {stage023[86]},
      {stage023[185]}
   );
   gpc1_1 gpc1_1_763(
      {stage023[87]},
      {stage023[186]}
   );
   gpc1_1 gpc1_1_764(
      {stage023[88]},
      {stage023[187]}
   );
   gpc1_1 gpc1_1_765(
      {stage023[89]},
      {stage023[188]}
   );
   gpc1_1 gpc1_1_766(
      {stage023[90]},
      {stage023[189]}
   );
   gpc1_1 gpc1_1_767(
      {stage023[91]},
      {stage023[190]}
   );
   gpc1_1 gpc1_1_768(
      {stage023[92]},
      {stage023[191]}
   );
   gpc1_1 gpc1_1_769(
      {stage023[93]},
      {stage023[192]}
   );
   gpc1_1 gpc1_1_770(
      {stage023[94]},
      {stage023[193]}
   );
   gpc1_1 gpc1_1_771(
      {stage023[95]},
      {stage023[194]}
   );
   gpc1_1 gpc1_1_772(
      {stage023[96]},
      {stage023[195]}
   );
   gpc1_1 gpc1_1_773(
      {stage023[97]},
      {stage023[196]}
   );
   gpc1_1 gpc1_1_774(
      {stage023[98]},
      {stage023[197]}
   );
   gpc1_1 gpc1_1_775(
      {stage023[99]},
      {stage023[198]}
   );
   gpc1_1 gpc1_1_776(
      {stage023[100]},
      {stage023[199]}
   );
   gpc1_1 gpc1_1_777(
      {stage023[101]},
      {stage023[200]}
   );
   gpc1_1 gpc1_1_778(
      {stage023[102]},
      {stage023[201]}
   );
   gpc1_1 gpc1_1_779(
      {stage023[103]},
      {stage023[202]}
   );
   gpc1_1 gpc1_1_780(
      {stage023[104]},
      {stage023[203]}
   );
   gpc1_1 gpc1_1_781(
      {stage023[105]},
      {stage023[204]}
   );
   gpc1_1 gpc1_1_782(
      {stage023[106]},
      {stage023[205]}
   );
   gpc1_1 gpc1_1_783(
      {stage023[107]},
      {stage023[206]}
   );
   gpc1_1 gpc1_1_784(
      {stage023[108]},
      {stage023[207]}
   );
   gpc1_1 gpc1_1_785(
      {stage023[109]},
      {stage023[208]}
   );
   gpc1_1 gpc1_1_786(
      {stage023[110]},
      {stage023[209]}
   );
   gpc1_1 gpc1_1_787(
      {stage023[111]},
      {stage023[210]}
   );
   gpc1_1 gpc1_1_788(
      {stage023[112]},
      {stage023[211]}
   );
   gpc1_1 gpc1_1_789(
      {stage023[113]},
      {stage023[212]}
   );
   gpc1_1 gpc1_1_790(
      {stage023[114]},
      {stage023[213]}
   );
   gpc1_1 gpc1_1_791(
      {stage023[115]},
      {stage023[214]}
   );
   gpc1_1 gpc1_1_792(
      {stage023[116]},
      {stage023[215]}
   );
   gpc1_1 gpc1_1_793(
      {stage023[117]},
      {stage023[216]}
   );
   gpc1_1 gpc1_1_794(
      {stage023[118]},
      {stage023[217]}
   );
   gpc1_1 gpc1_1_795(
      {stage023[119]},
      {stage023[218]}
   );
   gpc1_1 gpc1_1_796(
      {stage023[120]},
      {stage023[219]}
   );
   gpc1_1 gpc1_1_797(
      {stage023[121]},
      {stage023[220]}
   );
   gpc1_1 gpc1_1_798(
      {stage023[122]},
      {stage023[221]}
   );
   gpc1325_5 gpc1325_5_799(
      {stage023[123], stage023[124], stage023[125], stage023[126], stage023[127]},
      {stage024[60], stage024[61]},
      {stage025[0], stage025[1], stage025[2]},
      {stage026[0]},
      {stage027[128], stage026[138], stage025[148], stage024[158], stage023[222]}
   );
   gpc1_1 gpc1_1_800(
      {stage024[62]},
      {stage024[159]}
   );
   gpc1_1 gpc1_1_801(
      {stage024[63]},
      {stage024[160]}
   );
   gpc1_1 gpc1_1_802(
      {stage024[64]},
      {stage024[161]}
   );
   gpc1_1 gpc1_1_803(
      {stage024[65]},
      {stage024[162]}
   );
   gpc1_1 gpc1_1_804(
      {stage024[66]},
      {stage024[163]}
   );
   gpc1_1 gpc1_1_805(
      {stage024[67]},
      {stage024[164]}
   );
   gpc1_1 gpc1_1_806(
      {stage024[68]},
      {stage024[165]}
   );
   gpc1_1 gpc1_1_807(
      {stage024[69]},
      {stage024[166]}
   );
   gpc1_1 gpc1_1_808(
      {stage024[70]},
      {stage024[167]}
   );
   gpc1_1 gpc1_1_809(
      {stage024[71]},
      {stage024[168]}
   );
   gpc1_1 gpc1_1_810(
      {stage024[72]},
      {stage024[169]}
   );
   gpc1_1 gpc1_1_811(
      {stage024[73]},
      {stage024[170]}
   );
   gpc1_1 gpc1_1_812(
      {stage024[74]},
      {stage024[171]}
   );
   gpc1_1 gpc1_1_813(
      {stage024[75]},
      {stage024[172]}
   );
   gpc1_1 gpc1_1_814(
      {stage024[76]},
      {stage024[173]}
   );
   gpc1_1 gpc1_1_815(
      {stage024[77]},
      {stage024[174]}
   );
   gpc1_1 gpc1_1_816(
      {stage024[78]},
      {stage024[175]}
   );
   gpc1_1 gpc1_1_817(
      {stage024[79]},
      {stage024[176]}
   );
   gpc1_1 gpc1_1_818(
      {stage024[80]},
      {stage024[177]}
   );
   gpc1_1 gpc1_1_819(
      {stage024[81]},
      {stage024[178]}
   );
   gpc1_1 gpc1_1_820(
      {stage024[82]},
      {stage024[179]}
   );
   gpc606_5 gpc606_5_821(
      {stage024[83], stage024[84], stage024[85], stage024[86], stage024[87], stage024[88]},
      {stage026[1], stage026[2], stage026[3], stage026[4], stage026[5], stage026[6]},
      {stage028[128], stage027[129], stage026[139], stage025[149], stage024[180]}
   );
   gpc606_5 gpc606_5_822(
      {stage024[89], stage024[90], stage024[91], stage024[92], stage024[93], stage024[94]},
      {stage026[7], stage026[8], stage026[9], stage026[10], stage026[11], stage026[12]},
      {stage028[129], stage027[130], stage026[140], stage025[150], stage024[181]}
   );
   gpc606_5 gpc606_5_823(
      {stage024[95], stage024[96], stage024[97], stage024[98], stage024[99], stage024[100]},
      {stage026[13], stage026[14], stage026[15], stage026[16], stage026[17], stage026[18]},
      {stage028[130], stage027[131], stage026[141], stage025[151], stage024[182]}
   );
   gpc606_5 gpc606_5_824(
      {stage024[101], stage024[102], stage024[103], stage024[104], stage024[105], stage024[106]},
      {stage026[19], stage026[20], stage026[21], stage026[22], stage026[23], stage026[24]},
      {stage028[131], stage027[132], stage026[142], stage025[152], stage024[183]}
   );
   gpc606_5 gpc606_5_825(
      {stage024[107], stage024[108], stage024[109], stage024[110], stage024[111], stage024[112]},
      {stage026[25], stage026[26], stage026[27], stage026[28], stage026[29], stage026[30]},
      {stage028[132], stage027[133], stage026[143], stage025[153], stage024[184]}
   );
   gpc615_5 gpc615_5_826(
      {stage024[113], stage024[114], stage024[115], stage024[116], stage024[117]},
      {stage025[3]},
      {stage026[31], stage026[32], stage026[33], stage026[34], stage026[35], stage026[36]},
      {stage028[133], stage027[134], stage026[144], stage025[154], stage024[185]}
   );
   gpc615_5 gpc615_5_827(
      {stage024[118], stage024[119], stage024[120], stage024[121], stage024[122]},
      {stage025[4]},
      {stage026[37], stage026[38], stage026[39], stage026[40], stage026[41], stage026[42]},
      {stage028[134], stage027[135], stage026[145], stage025[155], stage024[186]}
   );
   gpc615_5 gpc615_5_828(
      {stage024[123], stage024[124], stage024[125], stage024[126], stage024[127]},
      {stage025[5]},
      {stage026[43], stage026[44], stage026[45], stage026[46], stage026[47], stage026[48]},
      {stage028[135], stage027[136], stage026[146], stage025[156], stage024[187]}
   );
   gpc1_1 gpc1_1_829(
      {stage025[6]},
      {stage025[157]}
   );
   gpc1_1 gpc1_1_830(
      {stage025[7]},
      {stage025[158]}
   );
   gpc1_1 gpc1_1_831(
      {stage025[8]},
      {stage025[159]}
   );
   gpc1_1 gpc1_1_832(
      {stage025[9]},
      {stage025[160]}
   );
   gpc1_1 gpc1_1_833(
      {stage025[10]},
      {stage025[161]}
   );
   gpc1_1 gpc1_1_834(
      {stage025[11]},
      {stage025[162]}
   );
   gpc1_1 gpc1_1_835(
      {stage025[12]},
      {stage025[163]}
   );
   gpc1_1 gpc1_1_836(
      {stage025[13]},
      {stage025[164]}
   );
   gpc1_1 gpc1_1_837(
      {stage025[14]},
      {stage025[165]}
   );
   gpc1_1 gpc1_1_838(
      {stage025[15]},
      {stage025[166]}
   );
   gpc1_1 gpc1_1_839(
      {stage025[16]},
      {stage025[167]}
   );
   gpc1_1 gpc1_1_840(
      {stage025[17]},
      {stage025[168]}
   );
   gpc1_1 gpc1_1_841(
      {stage025[18]},
      {stage025[169]}
   );
   gpc1_1 gpc1_1_842(
      {stage025[19]},
      {stage025[170]}
   );
   gpc1_1 gpc1_1_843(
      {stage025[20]},
      {stage025[171]}
   );
   gpc1_1 gpc1_1_844(
      {stage025[21]},
      {stage025[172]}
   );
   gpc1_1 gpc1_1_845(
      {stage025[22]},
      {stage025[173]}
   );
   gpc1_1 gpc1_1_846(
      {stage025[23]},
      {stage025[174]}
   );
   gpc1_1 gpc1_1_847(
      {stage025[24]},
      {stage025[175]}
   );
   gpc1_1 gpc1_1_848(
      {stage025[25]},
      {stage025[176]}
   );
   gpc1_1 gpc1_1_849(
      {stage025[26]},
      {stage025[177]}
   );
   gpc1_1 gpc1_1_850(
      {stage025[27]},
      {stage025[178]}
   );
   gpc1_1 gpc1_1_851(
      {stage025[28]},
      {stage025[179]}
   );
   gpc1_1 gpc1_1_852(
      {stage025[29]},
      {stage025[180]}
   );
   gpc1_1 gpc1_1_853(
      {stage025[30]},
      {stage025[181]}
   );
   gpc1_1 gpc1_1_854(
      {stage025[31]},
      {stage025[182]}
   );
   gpc1_1 gpc1_1_855(
      {stage025[32]},
      {stage025[183]}
   );
   gpc1_1 gpc1_1_856(
      {stage025[33]},
      {stage025[184]}
   );
   gpc1_1 gpc1_1_857(
      {stage025[34]},
      {stage025[185]}
   );
   gpc1_1 gpc1_1_858(
      {stage025[35]},
      {stage025[186]}
   );
   gpc1_1 gpc1_1_859(
      {stage025[36]},
      {stage025[187]}
   );
   gpc1_1 gpc1_1_860(
      {stage025[37]},
      {stage025[188]}
   );
   gpc1_1 gpc1_1_861(
      {stage025[38]},
      {stage025[189]}
   );
   gpc1_1 gpc1_1_862(
      {stage025[39]},
      {stage025[190]}
   );
   gpc1_1 gpc1_1_863(
      {stage025[40]},
      {stage025[191]}
   );
   gpc1_1 gpc1_1_864(
      {stage025[41]},
      {stage025[192]}
   );
   gpc1_1 gpc1_1_865(
      {stage025[42]},
      {stage025[193]}
   );
   gpc1_1 gpc1_1_866(
      {stage025[43]},
      {stage025[194]}
   );
   gpc1_1 gpc1_1_867(
      {stage025[44]},
      {stage025[195]}
   );
   gpc1_1 gpc1_1_868(
      {stage025[45]},
      {stage025[196]}
   );
   gpc1_1 gpc1_1_869(
      {stage025[46]},
      {stage025[197]}
   );
   gpc1_1 gpc1_1_870(
      {stage025[47]},
      {stage025[198]}
   );
   gpc1_1 gpc1_1_871(
      {stage025[48]},
      {stage025[199]}
   );
   gpc1_1 gpc1_1_872(
      {stage025[49]},
      {stage025[200]}
   );
   gpc1_1 gpc1_1_873(
      {stage025[50]},
      {stage025[201]}
   );
   gpc1_1 gpc1_1_874(
      {stage025[51]},
      {stage025[202]}
   );
   gpc1_1 gpc1_1_875(
      {stage025[52]},
      {stage025[203]}
   );
   gpc1_1 gpc1_1_876(
      {stage025[53]},
      {stage025[204]}
   );
   gpc1_1 gpc1_1_877(
      {stage025[54]},
      {stage025[205]}
   );
   gpc1_1 gpc1_1_878(
      {stage025[55]},
      {stage025[206]}
   );
   gpc623_5 gpc623_5_879(
      {stage025[56], stage025[57], stage025[58]},
      {stage026[49], stage026[50]},
      {stage027[0], stage027[1], stage027[2], stage027[3], stage027[4], stage027[5]},
      {stage029[128], stage028[136], stage027[137], stage026[147], stage025[207]}
   );
   gpc623_5 gpc623_5_880(
      {stage025[59], stage025[60], stage025[61]},
      {stage026[51], stage026[52]},
      {stage027[6], stage027[7], stage027[8], stage027[9], stage027[10], stage027[11]},
      {stage029[129], stage028[137], stage027[138], stage026[148], stage025[208]}
   );
   gpc623_5 gpc623_5_881(
      {stage025[62], stage025[63], stage025[64]},
      {stage026[53], stage026[54]},
      {stage027[12], stage027[13], stage027[14], stage027[15], stage027[16], stage027[17]},
      {stage029[130], stage028[138], stage027[139], stage026[149], stage025[209]}
   );
   gpc623_5 gpc623_5_882(
      {stage025[65], stage025[66], stage025[67]},
      {stage026[55], stage026[56]},
      {stage027[18], stage027[19], stage027[20], stage027[21], stage027[22], stage027[23]},
      {stage029[131], stage028[139], stage027[140], stage026[150], stage025[210]}
   );
   gpc623_5 gpc623_5_883(
      {stage025[68], stage025[69], stage025[70]},
      {stage026[57], stage026[58]},
      {stage027[24], stage027[25], stage027[26], stage027[27], stage027[28], stage027[29]},
      {stage029[132], stage028[140], stage027[141], stage026[151], stage025[211]}
   );
   gpc623_5 gpc623_5_884(
      {stage025[71], stage025[72], stage025[73]},
      {stage026[59], stage026[60]},
      {stage027[30], stage027[31], stage027[32], stage027[33], stage027[34], stage027[35]},
      {stage029[133], stage028[141], stage027[142], stage026[152], stage025[212]}
   );
   gpc623_5 gpc623_5_885(
      {stage025[74], stage025[75], stage025[76]},
      {stage026[61], stage026[62]},
      {stage027[36], stage027[37], stage027[38], stage027[39], stage027[40], stage027[41]},
      {stage029[134], stage028[142], stage027[143], stage026[153], stage025[213]}
   );
   gpc623_5 gpc623_5_886(
      {stage025[77], stage025[78], stage025[79]},
      {stage026[63], stage026[64]},
      {stage027[42], stage027[43], stage027[44], stage027[45], stage027[46], stage027[47]},
      {stage029[135], stage028[143], stage027[144], stage026[154], stage025[214]}
   );
   gpc623_5 gpc623_5_887(
      {stage025[80], stage025[81], stage025[82]},
      {stage026[65], stage026[66]},
      {stage027[48], stage027[49], stage027[50], stage027[51], stage027[52], stage027[53]},
      {stage029[136], stage028[144], stage027[145], stage026[155], stage025[215]}
   );
   gpc623_5 gpc623_5_888(
      {stage025[83], stage025[84], stage025[85]},
      {stage026[67], stage026[68]},
      {stage027[54], stage027[55], stage027[56], stage027[57], stage027[58], stage027[59]},
      {stage029[137], stage028[145], stage027[146], stage026[156], stage025[216]}
   );
   gpc606_5 gpc606_5_889(
      {stage025[86], stage025[87], stage025[88], stage025[89], stage025[90], stage025[91]},
      {stage027[60], stage027[61], stage027[62], stage027[63], stage027[64], stage027[65]},
      {stage029[138], stage028[146], stage027[147], stage026[157], stage025[217]}
   );
   gpc606_5 gpc606_5_890(
      {stage025[92], stage025[93], stage025[94], stage025[95], stage025[96], stage025[97]},
      {stage027[66], stage027[67], stage027[68], stage027[69], stage027[70], stage027[71]},
      {stage029[139], stage028[147], stage027[148], stage026[158], stage025[218]}
   );
   gpc606_5 gpc606_5_891(
      {stage025[98], stage025[99], stage025[100], stage025[101], stage025[102], stage025[103]},
      {stage027[72], stage027[73], stage027[74], stage027[75], stage027[76], stage027[77]},
      {stage029[140], stage028[148], stage027[149], stage026[159], stage025[219]}
   );
   gpc606_5 gpc606_5_892(
      {stage025[104], stage025[105], stage025[106], stage025[107], stage025[108], stage025[109]},
      {stage027[78], stage027[79], stage027[80], stage027[81], stage027[82], stage027[83]},
      {stage029[141], stage028[149], stage027[150], stage026[160], stage025[220]}
   );
   gpc606_5 gpc606_5_893(
      {stage025[110], stage025[111], stage025[112], stage025[113], stage025[114], stage025[115]},
      {stage027[84], stage027[85], stage027[86], stage027[87], stage027[88], stage027[89]},
      {stage029[142], stage028[150], stage027[151], stage026[161], stage025[221]}
   );
   gpc606_5 gpc606_5_894(
      {stage025[116], stage025[117], stage025[118], stage025[119], stage025[120], stage025[121]},
      {stage027[90], stage027[91], stage027[92], stage027[93], stage027[94], stage027[95]},
      {stage029[143], stage028[151], stage027[152], stage026[162], stage025[222]}
   );
   gpc606_5 gpc606_5_895(
      {stage025[122], stage025[123], stage025[124], stage025[125], stage025[126], stage025[127]},
      {stage027[96], stage027[97], stage027[98], stage027[99], stage027[100], stage027[101]},
      {stage029[144], stage028[152], stage027[153], stage026[163], stage025[223]}
   );
   gpc1_1 gpc1_1_896(
      {stage026[69]},
      {stage026[164]}
   );
   gpc1_1 gpc1_1_897(
      {stage026[70]},
      {stage026[165]}
   );
   gpc1_1 gpc1_1_898(
      {stage026[71]},
      {stage026[166]}
   );
   gpc1_1 gpc1_1_899(
      {stage026[72]},
      {stage026[167]}
   );
   gpc1_1 gpc1_1_900(
      {stage026[73]},
      {stage026[168]}
   );
   gpc1_1 gpc1_1_901(
      {stage026[74]},
      {stage026[169]}
   );
   gpc1_1 gpc1_1_902(
      {stage026[75]},
      {stage026[170]}
   );
   gpc1_1 gpc1_1_903(
      {stage026[76]},
      {stage026[171]}
   );
   gpc1_1 gpc1_1_904(
      {stage026[77]},
      {stage026[172]}
   );
   gpc1_1 gpc1_1_905(
      {stage026[78]},
      {stage026[173]}
   );
   gpc1_1 gpc1_1_906(
      {stage026[79]},
      {stage026[174]}
   );
   gpc1_1 gpc1_1_907(
      {stage026[80]},
      {stage026[175]}
   );
   gpc1_1 gpc1_1_908(
      {stage026[81]},
      {stage026[176]}
   );
   gpc1_1 gpc1_1_909(
      {stage026[82]},
      {stage026[177]}
   );
   gpc1_1 gpc1_1_910(
      {stage026[83]},
      {stage026[178]}
   );
   gpc1_1 gpc1_1_911(
      {stage026[84]},
      {stage026[179]}
   );
   gpc1_1 gpc1_1_912(
      {stage026[85]},
      {stage026[180]}
   );
   gpc1_1 gpc1_1_913(
      {stage026[86]},
      {stage026[181]}
   );
   gpc1_1 gpc1_1_914(
      {stage026[87]},
      {stage026[182]}
   );
   gpc615_5 gpc615_5_915(
      {stage026[88], stage026[89], stage026[90], stage026[91], stage026[92]},
      {stage027[102]},
      {stage028[0], stage028[1], stage028[2], stage028[3], stage028[4], stage028[5]},
      {stage030[128], stage029[145], stage028[153], stage027[154], stage026[183]}
   );
   gpc615_5 gpc615_5_916(
      {stage026[93], stage026[94], stage026[95], stage026[96], stage026[97]},
      {stage027[103]},
      {stage028[6], stage028[7], stage028[8], stage028[9], stage028[10], stage028[11]},
      {stage030[129], stage029[146], stage028[154], stage027[155], stage026[184]}
   );
   gpc615_5 gpc615_5_917(
      {stage026[98], stage026[99], stage026[100], stage026[101], stage026[102]},
      {stage027[104]},
      {stage028[12], stage028[13], stage028[14], stage028[15], stage028[16], stage028[17]},
      {stage030[130], stage029[147], stage028[155], stage027[156], stage026[185]}
   );
   gpc615_5 gpc615_5_918(
      {stage026[103], stage026[104], stage026[105], stage026[106], stage026[107]},
      {stage027[105]},
      {stage028[18], stage028[19], stage028[20], stage028[21], stage028[22], stage028[23]},
      {stage030[131], stage029[148], stage028[156], stage027[157], stage026[186]}
   );
   gpc615_5 gpc615_5_919(
      {stage026[108], stage026[109], stage026[110], stage026[111], stage026[112]},
      {stage027[106]},
      {stage028[24], stage028[25], stage028[26], stage028[27], stage028[28], stage028[29]},
      {stage030[132], stage029[149], stage028[157], stage027[158], stage026[187]}
   );
   gpc615_5 gpc615_5_920(
      {stage026[113], stage026[114], stage026[115], stage026[116], stage026[117]},
      {stage027[107]},
      {stage028[30], stage028[31], stage028[32], stage028[33], stage028[34], stage028[35]},
      {stage030[133], stage029[150], stage028[158], stage027[159], stage026[188]}
   );
   gpc615_5 gpc615_5_921(
      {stage026[118], stage026[119], stage026[120], stage026[121], stage026[122]},
      {stage027[108]},
      {stage028[36], stage028[37], stage028[38], stage028[39], stage028[40], stage028[41]},
      {stage030[134], stage029[151], stage028[159], stage027[160], stage026[189]}
   );
   gpc615_5 gpc615_5_922(
      {stage026[123], stage026[124], stage026[125], stage026[126], stage026[127]},
      {stage027[109]},
      {stage028[42], stage028[43], stage028[44], stage028[45], stage028[46], stage028[47]},
      {stage030[135], stage029[152], stage028[160], stage027[161], stage026[190]}
   );
   gpc1_1 gpc1_1_923(
      {stage027[110]},
      {stage027[162]}
   );
   gpc1_1 gpc1_1_924(
      {stage027[111]},
      {stage027[163]}
   );
   gpc1_1 gpc1_1_925(
      {stage027[112]},
      {stage027[164]}
   );
   gpc1_1 gpc1_1_926(
      {stage027[113]},
      {stage027[165]}
   );
   gpc1_1 gpc1_1_927(
      {stage027[114]},
      {stage027[166]}
   );
   gpc1_1 gpc1_1_928(
      {stage027[115]},
      {stage027[167]}
   );
   gpc1_1 gpc1_1_929(
      {stage027[116]},
      {stage027[168]}
   );
   gpc1_1 gpc1_1_930(
      {stage027[117]},
      {stage027[169]}
   );
   gpc1_1 gpc1_1_931(
      {stage027[118]},
      {stage027[170]}
   );
   gpc1_1 gpc1_1_932(
      {stage027[119]},
      {stage027[171]}
   );
   gpc1_1 gpc1_1_933(
      {stage027[120]},
      {stage027[172]}
   );
   gpc1_1 gpc1_1_934(
      {stage027[121]},
      {stage027[173]}
   );
   gpc1_1 gpc1_1_935(
      {stage027[122]},
      {stage027[174]}
   );
   gpc615_5 gpc615_5_936(
      {stage027[123], stage027[124], stage027[125], stage027[126], stage027[127]},
      {stage028[48]},
      {stage029[0], stage029[1], stage029[2], stage029[3], stage029[4], stage029[5]},
      {stage031[128], stage030[136], stage029[153], stage028[161], stage027[175]}
   );
   gpc1_1 gpc1_1_937(
      {stage028[49]},
      {stage028[162]}
   );
   gpc1_1 gpc1_1_938(
      {stage028[50]},
      {stage028[163]}
   );
   gpc1_1 gpc1_1_939(
      {stage028[51]},
      {stage028[164]}
   );
   gpc1_1 gpc1_1_940(
      {stage028[52]},
      {stage028[165]}
   );
   gpc1_1 gpc1_1_941(
      {stage028[53]},
      {stage028[166]}
   );
   gpc1_1 gpc1_1_942(
      {stage028[54]},
      {stage028[167]}
   );
   gpc606_5 gpc606_5_943(
      {stage028[55], stage028[56], stage028[57], stage028[58], stage028[59], stage028[60]},
      {stage030[0], stage030[1], stage030[2], stage030[3], stage030[4], stage030[5]},
      {stage032[128], stage031[129], stage030[137], stage029[154], stage028[168]}
   );
   gpc606_5 gpc606_5_944(
      {stage028[61], stage028[62], stage028[63], stage028[64], stage028[65], stage028[66]},
      {stage030[6], stage030[7], stage030[8], stage030[9], stage030[10], stage030[11]},
      {stage032[129], stage031[130], stage030[138], stage029[155], stage028[169]}
   );
   gpc606_5 gpc606_5_945(
      {stage028[67], stage028[68], stage028[69], stage028[70], stage028[71], stage028[72]},
      {stage030[12], stage030[13], stage030[14], stage030[15], stage030[16], stage030[17]},
      {stage032[130], stage031[131], stage030[139], stage029[156], stage028[170]}
   );
   gpc615_5 gpc615_5_946(
      {stage028[73], stage028[74], stage028[75], stage028[76], stage028[77]},
      {stage029[6]},
      {stage030[18], stage030[19], stage030[20], stage030[21], stage030[22], stage030[23]},
      {stage032[131], stage031[132], stage030[140], stage029[157], stage028[171]}
   );
   gpc615_5 gpc615_5_947(
      {stage028[78], stage028[79], stage028[80], stage028[81], stage028[82]},
      {stage029[7]},
      {stage030[24], stage030[25], stage030[26], stage030[27], stage030[28], stage030[29]},
      {stage032[132], stage031[133], stage030[141], stage029[158], stage028[172]}
   );
   gpc615_5 gpc615_5_948(
      {stage028[83], stage028[84], stage028[85], stage028[86], stage028[87]},
      {stage029[8]},
      {stage030[30], stage030[31], stage030[32], stage030[33], stage030[34], stage030[35]},
      {stage032[133], stage031[134], stage030[142], stage029[159], stage028[173]}
   );
   gpc615_5 gpc615_5_949(
      {stage028[88], stage028[89], stage028[90], stage028[91], stage028[92]},
      {stage029[9]},
      {stage030[36], stage030[37], stage030[38], stage030[39], stage030[40], stage030[41]},
      {stage032[134], stage031[135], stage030[143], stage029[160], stage028[174]}
   );
   gpc615_5 gpc615_5_950(
      {stage028[93], stage028[94], stage028[95], stage028[96], stage028[97]},
      {stage029[10]},
      {stage030[42], stage030[43], stage030[44], stage030[45], stage030[46], stage030[47]},
      {stage032[135], stage031[136], stage030[144], stage029[161], stage028[175]}
   );
   gpc615_5 gpc615_5_951(
      {stage028[98], stage028[99], stage028[100], stage028[101], stage028[102]},
      {stage029[11]},
      {stage030[48], stage030[49], stage030[50], stage030[51], stage030[52], stage030[53]},
      {stage032[136], stage031[137], stage030[145], stage029[162], stage028[176]}
   );
   gpc615_5 gpc615_5_952(
      {stage028[103], stage028[104], stage028[105], stage028[106], stage028[107]},
      {stage029[12]},
      {stage030[54], stage030[55], stage030[56], stage030[57], stage030[58], stage030[59]},
      {stage032[137], stage031[138], stage030[146], stage029[163], stage028[177]}
   );
   gpc615_5 gpc615_5_953(
      {stage028[108], stage028[109], stage028[110], stage028[111], stage028[112]},
      {stage029[13]},
      {stage030[60], stage030[61], stage030[62], stage030[63], stage030[64], stage030[65]},
      {stage032[138], stage031[139], stage030[147], stage029[164], stage028[178]}
   );
   gpc615_5 gpc615_5_954(
      {stage028[113], stage028[114], stage028[115], stage028[116], stage028[117]},
      {stage029[14]},
      {stage030[66], stage030[67], stage030[68], stage030[69], stage030[70], stage030[71]},
      {stage032[139], stage031[140], stage030[148], stage029[165], stage028[179]}
   );
   gpc615_5 gpc615_5_955(
      {stage028[118], stage028[119], stage028[120], stage028[121], stage028[122]},
      {stage029[15]},
      {stage030[72], stage030[73], stage030[74], stage030[75], stage030[76], stage030[77]},
      {stage032[140], stage031[141], stage030[149], stage029[166], stage028[180]}
   );
   gpc615_5 gpc615_5_956(
      {stage028[123], stage028[124], stage028[125], stage028[126], stage028[127]},
      {stage029[16]},
      {stage030[78], stage030[79], stage030[80], stage030[81], stage030[82], stage030[83]},
      {stage032[141], stage031[142], stage030[150], stage029[167], stage028[181]}
   );
   gpc1_1 gpc1_1_957(
      {stage029[17]},
      {stage029[168]}
   );
   gpc1_1 gpc1_1_958(
      {stage029[18]},
      {stage029[169]}
   );
   gpc1_1 gpc1_1_959(
      {stage029[19]},
      {stage029[170]}
   );
   gpc1_1 gpc1_1_960(
      {stage029[20]},
      {stage029[171]}
   );
   gpc1_1 gpc1_1_961(
      {stage029[21]},
      {stage029[172]}
   );
   gpc1_1 gpc1_1_962(
      {stage029[22]},
      {stage029[173]}
   );
   gpc1_1 gpc1_1_963(
      {stage029[23]},
      {stage029[174]}
   );
   gpc1_1 gpc1_1_964(
      {stage029[24]},
      {stage029[175]}
   );
   gpc1_1 gpc1_1_965(
      {stage029[25]},
      {stage029[176]}
   );
   gpc1_1 gpc1_1_966(
      {stage029[26]},
      {stage029[177]}
   );
   gpc1_1 gpc1_1_967(
      {stage029[27]},
      {stage029[178]}
   );
   gpc1_1 gpc1_1_968(
      {stage029[28]},
      {stage029[179]}
   );
   gpc1_1 gpc1_1_969(
      {stage029[29]},
      {stage029[180]}
   );
   gpc1_1 gpc1_1_970(
      {stage029[30]},
      {stage029[181]}
   );
   gpc1_1 gpc1_1_971(
      {stage029[31]},
      {stage029[182]}
   );
   gpc1_1 gpc1_1_972(
      {stage029[32]},
      {stage029[183]}
   );
   gpc1_1 gpc1_1_973(
      {stage029[33]},
      {stage029[184]}
   );
   gpc1_1 gpc1_1_974(
      {stage029[34]},
      {stage029[185]}
   );
   gpc1_1 gpc1_1_975(
      {stage029[35]},
      {stage029[186]}
   );
   gpc1_1 gpc1_1_976(
      {stage029[36]},
      {stage029[187]}
   );
   gpc1_1 gpc1_1_977(
      {stage029[37]},
      {stage029[188]}
   );
   gpc606_5 gpc606_5_978(
      {stage029[38], stage029[39], stage029[40], stage029[41], stage029[42], stage029[43]},
      {stage031[0], stage031[1], stage031[2], stage031[3], stage031[4], stage031[5]},
      {stage033[128], stage032[142], stage031[143], stage030[151], stage029[189]}
   );
   gpc606_5 gpc606_5_979(
      {stage029[44], stage029[45], stage029[46], stage029[47], stage029[48], stage029[49]},
      {stage031[6], stage031[7], stage031[8], stage031[9], stage031[10], stage031[11]},
      {stage033[129], stage032[143], stage031[144], stage030[152], stage029[190]}
   );
   gpc606_5 gpc606_5_980(
      {stage029[50], stage029[51], stage029[52], stage029[53], stage029[54], stage029[55]},
      {stage031[12], stage031[13], stage031[14], stage031[15], stage031[16], stage031[17]},
      {stage033[130], stage032[144], stage031[145], stage030[153], stage029[191]}
   );
   gpc606_5 gpc606_5_981(
      {stage029[56], stage029[57], stage029[58], stage029[59], stage029[60], stage029[61]},
      {stage031[18], stage031[19], stage031[20], stage031[21], stage031[22], stage031[23]},
      {stage033[131], stage032[145], stage031[146], stage030[154], stage029[192]}
   );
   gpc606_5 gpc606_5_982(
      {stage029[62], stage029[63], stage029[64], stage029[65], stage029[66], stage029[67]},
      {stage031[24], stage031[25], stage031[26], stage031[27], stage031[28], stage031[29]},
      {stage033[132], stage032[146], stage031[147], stage030[155], stage029[193]}
   );
   gpc606_5 gpc606_5_983(
      {stage029[68], stage029[69], stage029[70], stage029[71], stage029[72], stage029[73]},
      {stage031[30], stage031[31], stage031[32], stage031[33], stage031[34], stage031[35]},
      {stage033[133], stage032[147], stage031[148], stage030[156], stage029[194]}
   );
   gpc606_5 gpc606_5_984(
      {stage029[74], stage029[75], stage029[76], stage029[77], stage029[78], stage029[79]},
      {stage031[36], stage031[37], stage031[38], stage031[39], stage031[40], stage031[41]},
      {stage033[134], stage032[148], stage031[149], stage030[157], stage029[195]}
   );
   gpc606_5 gpc606_5_985(
      {stage029[80], stage029[81], stage029[82], stage029[83], stage029[84], stage029[85]},
      {stage031[42], stage031[43], stage031[44], stage031[45], stage031[46], stage031[47]},
      {stage033[135], stage032[149], stage031[150], stage030[158], stage029[196]}
   );
   gpc606_5 gpc606_5_986(
      {stage029[86], stage029[87], stage029[88], stage029[89], stage029[90], stage029[91]},
      {stage031[48], stage031[49], stage031[50], stage031[51], stage031[52], stage031[53]},
      {stage033[136], stage032[150], stage031[151], stage030[159], stage029[197]}
   );
   gpc606_5 gpc606_5_987(
      {stage029[92], stage029[93], stage029[94], stage029[95], stage029[96], stage029[97]},
      {stage031[54], stage031[55], stage031[56], stage031[57], stage031[58], stage031[59]},
      {stage033[137], stage032[151], stage031[152], stage030[160], stage029[198]}
   );
   gpc606_5 gpc606_5_988(
      {stage029[98], stage029[99], stage029[100], stage029[101], stage029[102], stage029[103]},
      {stage031[60], stage031[61], stage031[62], stage031[63], stage031[64], stage031[65]},
      {stage033[138], stage032[152], stage031[153], stage030[161], stage029[199]}
   );
   gpc606_5 gpc606_5_989(
      {stage029[104], stage029[105], stage029[106], stage029[107], stage029[108], stage029[109]},
      {stage031[66], stage031[67], stage031[68], stage031[69], stage031[70], stage031[71]},
      {stage033[139], stage032[153], stage031[154], stage030[162], stage029[200]}
   );
   gpc606_5 gpc606_5_990(
      {stage029[110], stage029[111], stage029[112], stage029[113], stage029[114], stage029[115]},
      {stage031[72], stage031[73], stage031[74], stage031[75], stage031[76], stage031[77]},
      {stage033[140], stage032[154], stage031[155], stage030[163], stage029[201]}
   );
   gpc606_5 gpc606_5_991(
      {stage029[116], stage029[117], stage029[118], stage029[119], stage029[120], stage029[121]},
      {stage031[78], stage031[79], stage031[80], stage031[81], stage031[82], stage031[83]},
      {stage033[141], stage032[155], stage031[156], stage030[164], stage029[202]}
   );
   gpc606_5 gpc606_5_992(
      {stage029[122], stage029[123], stage029[124], stage029[125], stage029[126], stage029[127]},
      {stage031[84], stage031[85], stage031[86], stage031[87], stage031[88], stage031[89]},
      {stage033[142], stage032[156], stage031[157], stage030[165], stage029[203]}
   );
   gpc1_1 gpc1_1_993(
      {stage030[84]},
      {stage030[166]}
   );
   gpc1_1 gpc1_1_994(
      {stage030[85]},
      {stage030[167]}
   );
   gpc1_1 gpc1_1_995(
      {stage030[86]},
      {stage030[168]}
   );
   gpc1_1 gpc1_1_996(
      {stage030[87]},
      {stage030[169]}
   );
   gpc1_1 gpc1_1_997(
      {stage030[88]},
      {stage030[170]}
   );
   gpc1_1 gpc1_1_998(
      {stage030[89]},
      {stage030[171]}
   );
   gpc1_1 gpc1_1_999(
      {stage030[90]},
      {stage030[172]}
   );
   gpc1_1 gpc1_1_1000(
      {stage030[91]},
      {stage030[173]}
   );
   gpc1_1 gpc1_1_1001(
      {stage030[92]},
      {stage030[174]}
   );
   gpc1_1 gpc1_1_1002(
      {stage030[93]},
      {stage030[175]}
   );
   gpc1_1 gpc1_1_1003(
      {stage030[94]},
      {stage030[176]}
   );
   gpc623_5 gpc623_5_1004(
      {stage030[95], stage030[96], stage030[97]},
      {stage031[90], stage031[91]},
      {stage032[0], stage032[1], stage032[2], stage032[3], stage032[4], stage032[5]},
      {stage034[128], stage033[143], stage032[157], stage031[158], stage030[177]}
   );
   gpc615_5 gpc615_5_1005(
      {stage030[98], stage030[99], stage030[100], stage030[101], stage030[102]},
      {stage031[92]},
      {stage032[6], stage032[7], stage032[8], stage032[9], stage032[10], stage032[11]},
      {stage034[129], stage033[144], stage032[158], stage031[159], stage030[178]}
   );
   gpc615_5 gpc615_5_1006(
      {stage030[103], stage030[104], stage030[105], stage030[106], stage030[107]},
      {stage031[93]},
      {stage032[12], stage032[13], stage032[14], stage032[15], stage032[16], stage032[17]},
      {stage034[130], stage033[145], stage032[159], stage031[160], stage030[179]}
   );
   gpc615_5 gpc615_5_1007(
      {stage030[108], stage030[109], stage030[110], stage030[111], stage030[112]},
      {stage031[94]},
      {stage032[18], stage032[19], stage032[20], stage032[21], stage032[22], stage032[23]},
      {stage034[131], stage033[146], stage032[160], stage031[161], stage030[180]}
   );
   gpc615_5 gpc615_5_1008(
      {stage030[113], stage030[114], stage030[115], stage030[116], stage030[117]},
      {stage031[95]},
      {stage032[24], stage032[25], stage032[26], stage032[27], stage032[28], stage032[29]},
      {stage034[132], stage033[147], stage032[161], stage031[162], stage030[181]}
   );
   gpc615_5 gpc615_5_1009(
      {stage030[118], stage030[119], stage030[120], stage030[121], stage030[122]},
      {stage031[96]},
      {stage032[30], stage032[31], stage032[32], stage032[33], stage032[34], stage032[35]},
      {stage034[133], stage033[148], stage032[162], stage031[163], stage030[182]}
   );
   gpc615_5 gpc615_5_1010(
      {stage030[123], stage030[124], stage030[125], stage030[126], stage030[127]},
      {stage031[97]},
      {stage032[36], stage032[37], stage032[38], stage032[39], stage032[40], stage032[41]},
      {stage034[134], stage033[149], stage032[163], stage031[164], stage030[183]}
   );
   gpc1_1 gpc1_1_1011(
      {stage031[98]},
      {stage031[165]}
   );
   gpc606_5 gpc606_5_1012(
      {stage031[99], stage031[100], stage031[101], stage031[102], stage031[103], stage031[104]},
      {stage033[0], stage033[1], stage033[2], stage033[3], stage033[4], stage033[5]},
      {stage035[128], stage034[135], stage033[150], stage032[164], stage031[166]}
   );
   gpc606_5 gpc606_5_1013(
      {stage031[105], stage031[106], stage031[107], stage031[108], stage031[109], stage031[110]},
      {stage033[6], stage033[7], stage033[8], stage033[9], stage033[10], stage033[11]},
      {stage035[129], stage034[136], stage033[151], stage032[165], stage031[167]}
   );
   gpc606_5 gpc606_5_1014(
      {stage031[111], stage031[112], stage031[113], stage031[114], stage031[115], stage031[116]},
      {stage033[12], stage033[13], stage033[14], stage033[15], stage033[16], stage033[17]},
      {stage035[130], stage034[137], stage033[152], stage032[166], stage031[168]}
   );
   gpc606_5 gpc606_5_1015(
      {stage031[117], stage031[118], stage031[119], stage031[120], stage031[121], stage031[122]},
      {stage033[18], stage033[19], stage033[20], stage033[21], stage033[22], stage033[23]},
      {stage035[131], stage034[138], stage033[153], stage032[167], stage031[169]}
   );
   gpc615_5 gpc615_5_1016(
      {stage031[123], stage031[124], stage031[125], stage031[126], stage031[127]},
      {stage032[42]},
      {stage033[24], stage033[25], stage033[26], stage033[27], stage033[28], stage033[29]},
      {stage035[132], stage034[139], stage033[154], stage032[168], stage031[170]}
   );
   gpc1_1 gpc1_1_1017(
      {stage032[43]},
      {stage032[169]}
   );
   gpc1_1 gpc1_1_1018(
      {stage032[44]},
      {stage032[170]}
   );
   gpc1_1 gpc1_1_1019(
      {stage032[45]},
      {stage032[171]}
   );
   gpc1_1 gpc1_1_1020(
      {stage032[46]},
      {stage032[172]}
   );
   gpc1_1 gpc1_1_1021(
      {stage032[47]},
      {stage032[173]}
   );
   gpc1_1 gpc1_1_1022(
      {stage032[48]},
      {stage032[174]}
   );
   gpc1_1 gpc1_1_1023(
      {stage032[49]},
      {stage032[175]}
   );
   gpc1_1 gpc1_1_1024(
      {stage032[50]},
      {stage032[176]}
   );
   gpc1_1 gpc1_1_1025(
      {stage032[51]},
      {stage032[177]}
   );
   gpc1_1 gpc1_1_1026(
      {stage032[52]},
      {stage032[178]}
   );
   gpc1_1 gpc1_1_1027(
      {stage032[53]},
      {stage032[179]}
   );
   gpc1_1 gpc1_1_1028(
      {stage032[54]},
      {stage032[180]}
   );
   gpc1_1 gpc1_1_1029(
      {stage032[55]},
      {stage032[181]}
   );
   gpc1_1 gpc1_1_1030(
      {stage032[56]},
      {stage032[182]}
   );
   gpc1_1 gpc1_1_1031(
      {stage032[57]},
      {stage032[183]}
   );
   gpc1_1 gpc1_1_1032(
      {stage032[58]},
      {stage032[184]}
   );
   gpc1_1 gpc1_1_1033(
      {stage032[59]},
      {stage032[185]}
   );
   gpc1_1 gpc1_1_1034(
      {stage032[60]},
      {stage032[186]}
   );
   gpc1_1 gpc1_1_1035(
      {stage032[61]},
      {stage032[187]}
   );
   gpc1_1 gpc1_1_1036(
      {stage032[62]},
      {stage032[188]}
   );
   gpc1_1 gpc1_1_1037(
      {stage032[63]},
      {stage032[189]}
   );
   gpc1_1 gpc1_1_1038(
      {stage032[64]},
      {stage032[190]}
   );
   gpc1_1 gpc1_1_1039(
      {stage032[65]},
      {stage032[191]}
   );
   gpc1_1 gpc1_1_1040(
      {stage032[66]},
      {stage032[192]}
   );
   gpc1_1 gpc1_1_1041(
      {stage032[67]},
      {stage032[193]}
   );
   gpc1_1 gpc1_1_1042(
      {stage032[68]},
      {stage032[194]}
   );
   gpc1_1 gpc1_1_1043(
      {stage032[69]},
      {stage032[195]}
   );
   gpc1_1 gpc1_1_1044(
      {stage032[70]},
      {stage032[196]}
   );
   gpc1_1 gpc1_1_1045(
      {stage032[71]},
      {stage032[197]}
   );
   gpc1_1 gpc1_1_1046(
      {stage032[72]},
      {stage032[198]}
   );
   gpc1_1 gpc1_1_1047(
      {stage032[73]},
      {stage032[199]}
   );
   gpc1_1 gpc1_1_1048(
      {stage032[74]},
      {stage032[200]}
   );
   gpc1_1 gpc1_1_1049(
      {stage032[75]},
      {stage032[201]}
   );
   gpc1_1 gpc1_1_1050(
      {stage032[76]},
      {stage032[202]}
   );
   gpc1_1 gpc1_1_1051(
      {stage032[77]},
      {stage032[203]}
   );
   gpc1_1 gpc1_1_1052(
      {stage032[78]},
      {stage032[204]}
   );
   gpc1_1 gpc1_1_1053(
      {stage032[79]},
      {stage032[205]}
   );
   gpc1_1 gpc1_1_1054(
      {stage032[80]},
      {stage032[206]}
   );
   gpc1_1 gpc1_1_1055(
      {stage032[81]},
      {stage032[207]}
   );
   gpc1_1 gpc1_1_1056(
      {stage032[82]},
      {stage032[208]}
   );
   gpc1_1 gpc1_1_1057(
      {stage032[83]},
      {stage032[209]}
   );
   gpc1_1 gpc1_1_1058(
      {stage032[84]},
      {stage032[210]}
   );
   gpc1_1 gpc1_1_1059(
      {stage032[85]},
      {stage032[211]}
   );
   gpc1_1 gpc1_1_1060(
      {stage032[86]},
      {stage032[212]}
   );
   gpc1_1 gpc1_1_1061(
      {stage032[87]},
      {stage032[213]}
   );
   gpc1_1 gpc1_1_1062(
      {stage032[88]},
      {stage032[214]}
   );
   gpc1_1 gpc1_1_1063(
      {stage032[89]},
      {stage032[215]}
   );
   gpc1_1 gpc1_1_1064(
      {stage032[90]},
      {stage032[216]}
   );
   gpc7_3 gpc7_3_1065(
      {stage032[91], stage032[92], stage032[93], stage032[94], stage032[95], stage032[96], stage032[97]},
      {stage034[140], stage033[155], stage032[217]}
   );
   gpc606_5 gpc606_5_1066(
      {stage032[98], stage032[99], stage032[100], stage032[101], stage032[102], stage032[103]},
      {stage034[0], stage034[1], stage034[2], stage034[3], stage034[4], stage034[5]},
      {stage036[128], stage035[133], stage034[141], stage033[156], stage032[218]}
   );
   gpc606_5 gpc606_5_1067(
      {stage032[104], stage032[105], stage032[106], stage032[107], stage032[108], stage032[109]},
      {stage034[6], stage034[7], stage034[8], stage034[9], stage034[10], stage034[11]},
      {stage036[129], stage035[134], stage034[142], stage033[157], stage032[219]}
   );
   gpc606_5 gpc606_5_1068(
      {stage032[110], stage032[111], stage032[112], stage032[113], stage032[114], stage032[115]},
      {stage034[12], stage034[13], stage034[14], stage034[15], stage034[16], stage034[17]},
      {stage036[130], stage035[135], stage034[143], stage033[158], stage032[220]}
   );
   gpc606_5 gpc606_5_1069(
      {stage032[116], stage032[117], stage032[118], stage032[119], stage032[120], stage032[121]},
      {stage034[18], stage034[19], stage034[20], stage034[21], stage034[22], stage034[23]},
      {stage036[131], stage035[136], stage034[144], stage033[159], stage032[221]}
   );
   gpc606_5 gpc606_5_1070(
      {stage032[122], stage032[123], stage032[124], stage032[125], stage032[126], stage032[127]},
      {stage034[24], stage034[25], stage034[26], stage034[27], stage034[28], stage034[29]},
      {stage036[132], stage035[137], stage034[145], stage033[160], stage032[222]}
   );
   gpc1_1 gpc1_1_1071(
      {stage033[30]},
      {stage033[161]}
   );
   gpc1_1 gpc1_1_1072(
      {stage033[31]},
      {stage033[162]}
   );
   gpc1_1 gpc1_1_1073(
      {stage033[32]},
      {stage033[163]}
   );
   gpc1_1 gpc1_1_1074(
      {stage033[33]},
      {stage033[164]}
   );
   gpc1_1 gpc1_1_1075(
      {stage033[34]},
      {stage033[165]}
   );
   gpc1_1 gpc1_1_1076(
      {stage033[35]},
      {stage033[166]}
   );
   gpc1_1 gpc1_1_1077(
      {stage033[36]},
      {stage033[167]}
   );
   gpc1_1 gpc1_1_1078(
      {stage033[37]},
      {stage033[168]}
   );
   gpc1_1 gpc1_1_1079(
      {stage033[38]},
      {stage033[169]}
   );
   gpc1_1 gpc1_1_1080(
      {stage033[39]},
      {stage033[170]}
   );
   gpc1_1 gpc1_1_1081(
      {stage033[40]},
      {stage033[171]}
   );
   gpc1_1 gpc1_1_1082(
      {stage033[41]},
      {stage033[172]}
   );
   gpc1_1 gpc1_1_1083(
      {stage033[42]},
      {stage033[173]}
   );
   gpc1_1 gpc1_1_1084(
      {stage033[43]},
      {stage033[174]}
   );
   gpc1_1 gpc1_1_1085(
      {stage033[44]},
      {stage033[175]}
   );
   gpc1_1 gpc1_1_1086(
      {stage033[45]},
      {stage033[176]}
   );
   gpc1_1 gpc1_1_1087(
      {stage033[46]},
      {stage033[177]}
   );
   gpc1_1 gpc1_1_1088(
      {stage033[47]},
      {stage033[178]}
   );
   gpc1_1 gpc1_1_1089(
      {stage033[48]},
      {stage033[179]}
   );
   gpc1_1 gpc1_1_1090(
      {stage033[49]},
      {stage033[180]}
   );
   gpc1_1 gpc1_1_1091(
      {stage033[50]},
      {stage033[181]}
   );
   gpc1_1 gpc1_1_1092(
      {stage033[51]},
      {stage033[182]}
   );
   gpc1_1 gpc1_1_1093(
      {stage033[52]},
      {stage033[183]}
   );
   gpc1_1 gpc1_1_1094(
      {stage033[53]},
      {stage033[184]}
   );
   gpc1_1 gpc1_1_1095(
      {stage033[54]},
      {stage033[185]}
   );
   gpc1_1 gpc1_1_1096(
      {stage033[55]},
      {stage033[186]}
   );
   gpc1_1 gpc1_1_1097(
      {stage033[56]},
      {stage033[187]}
   );
   gpc1_1 gpc1_1_1098(
      {stage033[57]},
      {stage033[188]}
   );
   gpc1_1 gpc1_1_1099(
      {stage033[58]},
      {stage033[189]}
   );
   gpc1_1 gpc1_1_1100(
      {stage033[59]},
      {stage033[190]}
   );
   gpc1_1 gpc1_1_1101(
      {stage033[60]},
      {stage033[191]}
   );
   gpc1_1 gpc1_1_1102(
      {stage033[61]},
      {stage033[192]}
   );
   gpc1_1 gpc1_1_1103(
      {stage033[62]},
      {stage033[193]}
   );
   gpc1_1 gpc1_1_1104(
      {stage033[63]},
      {stage033[194]}
   );
   gpc1_1 gpc1_1_1105(
      {stage033[64]},
      {stage033[195]}
   );
   gpc1_1 gpc1_1_1106(
      {stage033[65]},
      {stage033[196]}
   );
   gpc1_1 gpc1_1_1107(
      {stage033[66]},
      {stage033[197]}
   );
   gpc1_1 gpc1_1_1108(
      {stage033[67]},
      {stage033[198]}
   );
   gpc1_1 gpc1_1_1109(
      {stage033[68]},
      {stage033[199]}
   );
   gpc1_1 gpc1_1_1110(
      {stage033[69]},
      {stage033[200]}
   );
   gpc1_1 gpc1_1_1111(
      {stage033[70]},
      {stage033[201]}
   );
   gpc1_1 gpc1_1_1112(
      {stage033[71]},
      {stage033[202]}
   );
   gpc1_1 gpc1_1_1113(
      {stage033[72]},
      {stage033[203]}
   );
   gpc1_1 gpc1_1_1114(
      {stage033[73]},
      {stage033[204]}
   );
   gpc1_1 gpc1_1_1115(
      {stage033[74]},
      {stage033[205]}
   );
   gpc1_1 gpc1_1_1116(
      {stage033[75]},
      {stage033[206]}
   );
   gpc606_5 gpc606_5_1117(
      {stage033[76], stage033[77], stage033[78], stage033[79], stage033[80], stage033[81]},
      {stage035[0], stage035[1], stage035[2], stage035[3], stage035[4], stage035[5]},
      {stage037[128], stage036[133], stage035[138], stage034[146], stage033[207]}
   );
   gpc606_5 gpc606_5_1118(
      {stage033[82], stage033[83], stage033[84], stage033[85], stage033[86], stage033[87]},
      {stage035[6], stage035[7], stage035[8], stage035[9], stage035[10], stage035[11]},
      {stage037[129], stage036[134], stage035[139], stage034[147], stage033[208]}
   );
   gpc606_5 gpc606_5_1119(
      {stage033[88], stage033[89], stage033[90], stage033[91], stage033[92], stage033[93]},
      {stage035[12], stage035[13], stage035[14], stage035[15], stage035[16], stage035[17]},
      {stage037[130], stage036[135], stage035[140], stage034[148], stage033[209]}
   );
   gpc606_5 gpc606_5_1120(
      {stage033[94], stage033[95], stage033[96], stage033[97], stage033[98], stage033[99]},
      {stage035[18], stage035[19], stage035[20], stage035[21], stage035[22], stage035[23]},
      {stage037[131], stage036[136], stage035[141], stage034[149], stage033[210]}
   );
   gpc606_5 gpc606_5_1121(
      {stage033[100], stage033[101], stage033[102], stage033[103], stage033[104], stage033[105]},
      {stage035[24], stage035[25], stage035[26], stage035[27], stage035[28], stage035[29]},
      {stage037[132], stage036[137], stage035[142], stage034[150], stage033[211]}
   );
   gpc606_5 gpc606_5_1122(
      {stage033[106], stage033[107], stage033[108], stage033[109], stage033[110], stage033[111]},
      {stage035[30], stage035[31], stage035[32], stage035[33], stage035[34], stage035[35]},
      {stage037[133], stage036[138], stage035[143], stage034[151], stage033[212]}
   );
   gpc606_5 gpc606_5_1123(
      {stage033[112], stage033[113], stage033[114], stage033[115], stage033[116], stage033[117]},
      {stage035[36], stage035[37], stage035[38], stage035[39], stage035[40], stage035[41]},
      {stage037[134], stage036[139], stage035[144], stage034[152], stage033[213]}
   );
   gpc615_5 gpc615_5_1124(
      {stage033[118], stage033[119], stage033[120], stage033[121], stage033[122]},
      {stage034[30]},
      {stage035[42], stage035[43], stage035[44], stage035[45], stage035[46], stage035[47]},
      {stage037[135], stage036[140], stage035[145], stage034[153], stage033[214]}
   );
   gpc615_5 gpc615_5_1125(
      {stage033[123], stage033[124], stage033[125], stage033[126], stage033[127]},
      {stage034[31]},
      {stage035[48], stage035[49], stage035[50], stage035[51], stage035[52], stage035[53]},
      {stage037[136], stage036[141], stage035[146], stage034[154], stage033[215]}
   );
   gpc1_1 gpc1_1_1126(
      {stage034[32]},
      {stage034[155]}
   );
   gpc1_1 gpc1_1_1127(
      {stage034[33]},
      {stage034[156]}
   );
   gpc1_1 gpc1_1_1128(
      {stage034[34]},
      {stage034[157]}
   );
   gpc1_1 gpc1_1_1129(
      {stage034[35]},
      {stage034[158]}
   );
   gpc1_1 gpc1_1_1130(
      {stage034[36]},
      {stage034[159]}
   );
   gpc1_1 gpc1_1_1131(
      {stage034[37]},
      {stage034[160]}
   );
   gpc1_1 gpc1_1_1132(
      {stage034[38]},
      {stage034[161]}
   );
   gpc1_1 gpc1_1_1133(
      {stage034[39]},
      {stage034[162]}
   );
   gpc1_1 gpc1_1_1134(
      {stage034[40]},
      {stage034[163]}
   );
   gpc1_1 gpc1_1_1135(
      {stage034[41]},
      {stage034[164]}
   );
   gpc1_1 gpc1_1_1136(
      {stage034[42]},
      {stage034[165]}
   );
   gpc1_1 gpc1_1_1137(
      {stage034[43]},
      {stage034[166]}
   );
   gpc1_1 gpc1_1_1138(
      {stage034[44]},
      {stage034[167]}
   );
   gpc1_1 gpc1_1_1139(
      {stage034[45]},
      {stage034[168]}
   );
   gpc1_1 gpc1_1_1140(
      {stage034[46]},
      {stage034[169]}
   );
   gpc1_1 gpc1_1_1141(
      {stage034[47]},
      {stage034[170]}
   );
   gpc1_1 gpc1_1_1142(
      {stage034[48]},
      {stage034[171]}
   );
   gpc1_1 gpc1_1_1143(
      {stage034[49]},
      {stage034[172]}
   );
   gpc1_1 gpc1_1_1144(
      {stage034[50]},
      {stage034[173]}
   );
   gpc1_1 gpc1_1_1145(
      {stage034[51]},
      {stage034[174]}
   );
   gpc1_1 gpc1_1_1146(
      {stage034[52]},
      {stage034[175]}
   );
   gpc1_1 gpc1_1_1147(
      {stage034[53]},
      {stage034[176]}
   );
   gpc1_1 gpc1_1_1148(
      {stage034[54]},
      {stage034[177]}
   );
   gpc1_1 gpc1_1_1149(
      {stage034[55]},
      {stage034[178]}
   );
   gpc1_1 gpc1_1_1150(
      {stage034[56]},
      {stage034[179]}
   );
   gpc1_1 gpc1_1_1151(
      {stage034[57]},
      {stage034[180]}
   );
   gpc1_1 gpc1_1_1152(
      {stage034[58]},
      {stage034[181]}
   );
   gpc1_1 gpc1_1_1153(
      {stage034[59]},
      {stage034[182]}
   );
   gpc1_1 gpc1_1_1154(
      {stage034[60]},
      {stage034[183]}
   );
   gpc1_1 gpc1_1_1155(
      {stage034[61]},
      {stage034[184]}
   );
   gpc1_1 gpc1_1_1156(
      {stage034[62]},
      {stage034[185]}
   );
   gpc1_1 gpc1_1_1157(
      {stage034[63]},
      {stage034[186]}
   );
   gpc1_1 gpc1_1_1158(
      {stage034[64]},
      {stage034[187]}
   );
   gpc1_1 gpc1_1_1159(
      {stage034[65]},
      {stage034[188]}
   );
   gpc1_1 gpc1_1_1160(
      {stage034[66]},
      {stage034[189]}
   );
   gpc1_1 gpc1_1_1161(
      {stage034[67]},
      {stage034[190]}
   );
   gpc1_1 gpc1_1_1162(
      {stage034[68]},
      {stage034[191]}
   );
   gpc1_1 gpc1_1_1163(
      {stage034[69]},
      {stage034[192]}
   );
   gpc1_1 gpc1_1_1164(
      {stage034[70]},
      {stage034[193]}
   );
   gpc1_1 gpc1_1_1165(
      {stage034[71]},
      {stage034[194]}
   );
   gpc1_1 gpc1_1_1166(
      {stage034[72]},
      {stage034[195]}
   );
   gpc1_1 gpc1_1_1167(
      {stage034[73]},
      {stage034[196]}
   );
   gpc1_1 gpc1_1_1168(
      {stage034[74]},
      {stage034[197]}
   );
   gpc1_1 gpc1_1_1169(
      {stage034[75]},
      {stage034[198]}
   );
   gpc1_1 gpc1_1_1170(
      {stage034[76]},
      {stage034[199]}
   );
   gpc1_1 gpc1_1_1171(
      {stage034[77]},
      {stage034[200]}
   );
   gpc615_5 gpc615_5_1172(
      {stage034[78], stage034[79], stage034[80], stage034[81], stage034[82]},
      {stage035[54]},
      {stage036[0], stage036[1], stage036[2], stage036[3], stage036[4], stage036[5]},
      {stage038[128], stage037[137], stage036[142], stage035[147], stage034[201]}
   );
   gpc615_5 gpc615_5_1173(
      {stage034[83], stage034[84], stage034[85], stage034[86], stage034[87]},
      {stage035[55]},
      {stage036[6], stage036[7], stage036[8], stage036[9], stage036[10], stage036[11]},
      {stage038[129], stage037[138], stage036[143], stage035[148], stage034[202]}
   );
   gpc615_5 gpc615_5_1174(
      {stage034[88], stage034[89], stage034[90], stage034[91], stage034[92]},
      {stage035[56]},
      {stage036[12], stage036[13], stage036[14], stage036[15], stage036[16], stage036[17]},
      {stage038[130], stage037[139], stage036[144], stage035[149], stage034[203]}
   );
   gpc615_5 gpc615_5_1175(
      {stage034[93], stage034[94], stage034[95], stage034[96], stage034[97]},
      {stage035[57]},
      {stage036[18], stage036[19], stage036[20], stage036[21], stage036[22], stage036[23]},
      {stage038[131], stage037[140], stage036[145], stage035[150], stage034[204]}
   );
   gpc615_5 gpc615_5_1176(
      {stage034[98], stage034[99], stage034[100], stage034[101], stage034[102]},
      {stage035[58]},
      {stage036[24], stage036[25], stage036[26], stage036[27], stage036[28], stage036[29]},
      {stage038[132], stage037[141], stage036[146], stage035[151], stage034[205]}
   );
   gpc615_5 gpc615_5_1177(
      {stage034[103], stage034[104], stage034[105], stage034[106], stage034[107]},
      {stage035[59]},
      {stage036[30], stage036[31], stage036[32], stage036[33], stage036[34], stage036[35]},
      {stage038[133], stage037[142], stage036[147], stage035[152], stage034[206]}
   );
   gpc615_5 gpc615_5_1178(
      {stage034[108], stage034[109], stage034[110], stage034[111], stage034[112]},
      {stage035[60]},
      {stage036[36], stage036[37], stage036[38], stage036[39], stage036[40], stage036[41]},
      {stage038[134], stage037[143], stage036[148], stage035[153], stage034[207]}
   );
   gpc615_5 gpc615_5_1179(
      {stage034[113], stage034[114], stage034[115], stage034[116], stage034[117]},
      {stage035[61]},
      {stage036[42], stage036[43], stage036[44], stage036[45], stage036[46], stage036[47]},
      {stage038[135], stage037[144], stage036[149], stage035[154], stage034[208]}
   );
   gpc1415_5 gpc1415_5_1180(
      {stage034[118], stage034[119], stage034[120], stage034[121], stage034[122]},
      {stage035[62]},
      {stage036[48], stage036[49], stage036[50], stage036[51]},
      {stage037[0]},
      {stage038[136], stage037[145], stage036[150], stage035[155], stage034[209]}
   );
   gpc1415_5 gpc1415_5_1181(
      {stage034[123], stage034[124], stage034[125], stage034[126], stage034[127]},
      {stage035[63]},
      {stage036[52], stage036[53], stage036[54], stage036[55]},
      {stage037[1]},
      {stage038[137], stage037[146], stage036[151], stage035[156], stage034[210]}
   );
   gpc1_1 gpc1_1_1182(
      {stage035[64]},
      {stage035[157]}
   );
   gpc1_1 gpc1_1_1183(
      {stage035[65]},
      {stage035[158]}
   );
   gpc1_1 gpc1_1_1184(
      {stage035[66]},
      {stage035[159]}
   );
   gpc1_1 gpc1_1_1185(
      {stage035[67]},
      {stage035[160]}
   );
   gpc1_1 gpc1_1_1186(
      {stage035[68]},
      {stage035[161]}
   );
   gpc1_1 gpc1_1_1187(
      {stage035[69]},
      {stage035[162]}
   );
   gpc1_1 gpc1_1_1188(
      {stage035[70]},
      {stage035[163]}
   );
   gpc1_1 gpc1_1_1189(
      {stage035[71]},
      {stage035[164]}
   );
   gpc1_1 gpc1_1_1190(
      {stage035[72]},
      {stage035[165]}
   );
   gpc1_1 gpc1_1_1191(
      {stage035[73]},
      {stage035[166]}
   );
   gpc1_1 gpc1_1_1192(
      {stage035[74]},
      {stage035[167]}
   );
   gpc1_1 gpc1_1_1193(
      {stage035[75]},
      {stage035[168]}
   );
   gpc1_1 gpc1_1_1194(
      {stage035[76]},
      {stage035[169]}
   );
   gpc1_1 gpc1_1_1195(
      {stage035[77]},
      {stage035[170]}
   );
   gpc1_1 gpc1_1_1196(
      {stage035[78]},
      {stage035[171]}
   );
   gpc1_1 gpc1_1_1197(
      {stage035[79]},
      {stage035[172]}
   );
   gpc1_1 gpc1_1_1198(
      {stage035[80]},
      {stage035[173]}
   );
   gpc1_1 gpc1_1_1199(
      {stage035[81]},
      {stage035[174]}
   );
   gpc1_1 gpc1_1_1200(
      {stage035[82]},
      {stage035[175]}
   );
   gpc1_1 gpc1_1_1201(
      {stage035[83]},
      {stage035[176]}
   );
   gpc1_1 gpc1_1_1202(
      {stage035[84]},
      {stage035[177]}
   );
   gpc1_1 gpc1_1_1203(
      {stage035[85]},
      {stage035[178]}
   );
   gpc1_1 gpc1_1_1204(
      {stage035[86]},
      {stage035[179]}
   );
   gpc1_1 gpc1_1_1205(
      {stage035[87]},
      {stage035[180]}
   );
   gpc1_1 gpc1_1_1206(
      {stage035[88]},
      {stage035[181]}
   );
   gpc1_1 gpc1_1_1207(
      {stage035[89]},
      {stage035[182]}
   );
   gpc1_1 gpc1_1_1208(
      {stage035[90]},
      {stage035[183]}
   );
   gpc1_1 gpc1_1_1209(
      {stage035[91]},
      {stage035[184]}
   );
   gpc1_1 gpc1_1_1210(
      {stage035[92]},
      {stage035[185]}
   );
   gpc1_1 gpc1_1_1211(
      {stage035[93]},
      {stage035[186]}
   );
   gpc1_1 gpc1_1_1212(
      {stage035[94]},
      {stage035[187]}
   );
   gpc1_1 gpc1_1_1213(
      {stage035[95]},
      {stage035[188]}
   );
   gpc1_1 gpc1_1_1214(
      {stage035[96]},
      {stage035[189]}
   );
   gpc1_1 gpc1_1_1215(
      {stage035[97]},
      {stage035[190]}
   );
   gpc1_1 gpc1_1_1216(
      {stage035[98]},
      {stage035[191]}
   );
   gpc1_1 gpc1_1_1217(
      {stage035[99]},
      {stage035[192]}
   );
   gpc1_1 gpc1_1_1218(
      {stage035[100]},
      {stage035[193]}
   );
   gpc1_1 gpc1_1_1219(
      {stage035[101]},
      {stage035[194]}
   );
   gpc1_1 gpc1_1_1220(
      {stage035[102]},
      {stage035[195]}
   );
   gpc1_1 gpc1_1_1221(
      {stage035[103]},
      {stage035[196]}
   );
   gpc1_1 gpc1_1_1222(
      {stage035[104]},
      {stage035[197]}
   );
   gpc1_1 gpc1_1_1223(
      {stage035[105]},
      {stage035[198]}
   );
   gpc1_1 gpc1_1_1224(
      {stage035[106]},
      {stage035[199]}
   );
   gpc1_1 gpc1_1_1225(
      {stage035[107]},
      {stage035[200]}
   );
   gpc1_1 gpc1_1_1226(
      {stage035[108]},
      {stage035[201]}
   );
   gpc1_1 gpc1_1_1227(
      {stage035[109]},
      {stage035[202]}
   );
   gpc1_1 gpc1_1_1228(
      {stage035[110]},
      {stage035[203]}
   );
   gpc1_1 gpc1_1_1229(
      {stage035[111]},
      {stage035[204]}
   );
   gpc1_1 gpc1_1_1230(
      {stage035[112]},
      {stage035[205]}
   );
   gpc615_5 gpc615_5_1231(
      {stage035[113], stage035[114], stage035[115], stage035[116], stage035[117]},
      {stage036[56]},
      {stage037[2], stage037[3], stage037[4], stage037[5], stage037[6], stage037[7]},
      {stage039[128], stage038[138], stage037[147], stage036[152], stage035[206]}
   );
   gpc615_5 gpc615_5_1232(
      {stage035[118], stage035[119], stage035[120], stage035[121], stage035[122]},
      {stage036[57]},
      {stage037[8], stage037[9], stage037[10], stage037[11], stage037[12], stage037[13]},
      {stage039[129], stage038[139], stage037[148], stage036[153], stage035[207]}
   );
   gpc2135_5 gpc2135_5_1233(
      {stage035[123], stage035[124], stage035[125], stage035[126], stage035[127]},
      {stage036[58], stage036[59], stage036[60]},
      {stage037[14]},
      {stage038[0], stage038[1]},
      {stage039[130], stage038[140], stage037[149], stage036[154], stage035[208]}
   );
   gpc1_1 gpc1_1_1234(
      {stage036[61]},
      {stage036[155]}
   );
   gpc1_1 gpc1_1_1235(
      {stage036[62]},
      {stage036[156]}
   );
   gpc1_1 gpc1_1_1236(
      {stage036[63]},
      {stage036[157]}
   );
   gpc1_1 gpc1_1_1237(
      {stage036[64]},
      {stage036[158]}
   );
   gpc1_1 gpc1_1_1238(
      {stage036[65]},
      {stage036[159]}
   );
   gpc1_1 gpc1_1_1239(
      {stage036[66]},
      {stage036[160]}
   );
   gpc1_1 gpc1_1_1240(
      {stage036[67]},
      {stage036[161]}
   );
   gpc1_1 gpc1_1_1241(
      {stage036[68]},
      {stage036[162]}
   );
   gpc606_5 gpc606_5_1242(
      {stage036[69], stage036[70], stage036[71], stage036[72], stage036[73], stage036[74]},
      {stage038[2], stage038[3], stage038[4], stage038[5], stage038[6], stage038[7]},
      {stage040[128], stage039[131], stage038[141], stage037[150], stage036[163]}
   );
   gpc606_5 gpc606_5_1243(
      {stage036[75], stage036[76], stage036[77], stage036[78], stage036[79], stage036[80]},
      {stage038[8], stage038[9], stage038[10], stage038[11], stage038[12], stage038[13]},
      {stage040[129], stage039[132], stage038[142], stage037[151], stage036[164]}
   );
   gpc606_5 gpc606_5_1244(
      {stage036[81], stage036[82], stage036[83], stage036[84], stage036[85], stage036[86]},
      {stage038[14], stage038[15], stage038[16], stage038[17], stage038[18], stage038[19]},
      {stage040[130], stage039[133], stage038[143], stage037[152], stage036[165]}
   );
   gpc606_5 gpc606_5_1245(
      {stage036[87], stage036[88], stage036[89], stage036[90], stage036[91], stage036[92]},
      {stage038[20], stage038[21], stage038[22], stage038[23], stage038[24], stage038[25]},
      {stage040[131], stage039[134], stage038[144], stage037[153], stage036[166]}
   );
   gpc606_5 gpc606_5_1246(
      {stage036[93], stage036[94], stage036[95], stage036[96], stage036[97], stage036[98]},
      {stage038[26], stage038[27], stage038[28], stage038[29], stage038[30], stage038[31]},
      {stage040[132], stage039[135], stage038[145], stage037[154], stage036[167]}
   );
   gpc606_5 gpc606_5_1247(
      {stage036[99], stage036[100], stage036[101], stage036[102], stage036[103], stage036[104]},
      {stage038[32], stage038[33], stage038[34], stage038[35], stage038[36], stage038[37]},
      {stage040[133], stage039[136], stage038[146], stage037[155], stage036[168]}
   );
   gpc606_5 gpc606_5_1248(
      {stage036[105], stage036[106], stage036[107], stage036[108], stage036[109], stage036[110]},
      {stage038[38], stage038[39], stage038[40], stage038[41], stage038[42], stage038[43]},
      {stage040[134], stage039[137], stage038[147], stage037[156], stage036[169]}
   );
   gpc606_5 gpc606_5_1249(
      {stage036[111], stage036[112], stage036[113], stage036[114], stage036[115], stage036[116]},
      {stage038[44], stage038[45], stage038[46], stage038[47], stage038[48], stage038[49]},
      {stage040[135], stage039[138], stage038[148], stage037[157], stage036[170]}
   );
   gpc606_5 gpc606_5_1250(
      {stage036[117], stage036[118], stage036[119], stage036[120], stage036[121], stage036[122]},
      {stage038[50], stage038[51], stage038[52], stage038[53], stage038[54], stage038[55]},
      {stage040[136], stage039[139], stage038[149], stage037[158], stage036[171]}
   );
   gpc615_5 gpc615_5_1251(
      {stage036[123], stage036[124], stage036[125], stage036[126], stage036[127]},
      {stage037[15]},
      {stage038[56], stage038[57], stage038[58], stage038[59], stage038[60], stage038[61]},
      {stage040[137], stage039[140], stage038[150], stage037[159], stage036[172]}
   );
   gpc1_1 gpc1_1_1252(
      {stage037[16]},
      {stage037[160]}
   );
   gpc1_1 gpc1_1_1253(
      {stage037[17]},
      {stage037[161]}
   );
   gpc1_1 gpc1_1_1254(
      {stage037[18]},
      {stage037[162]}
   );
   gpc1_1 gpc1_1_1255(
      {stage037[19]},
      {stage037[163]}
   );
   gpc1_1 gpc1_1_1256(
      {stage037[20]},
      {stage037[164]}
   );
   gpc1_1 gpc1_1_1257(
      {stage037[21]},
      {stage037[165]}
   );
   gpc1_1 gpc1_1_1258(
      {stage037[22]},
      {stage037[166]}
   );
   gpc1_1 gpc1_1_1259(
      {stage037[23]},
      {stage037[167]}
   );
   gpc1_1 gpc1_1_1260(
      {stage037[24]},
      {stage037[168]}
   );
   gpc1_1 gpc1_1_1261(
      {stage037[25]},
      {stage037[169]}
   );
   gpc1_1 gpc1_1_1262(
      {stage037[26]},
      {stage037[170]}
   );
   gpc1_1 gpc1_1_1263(
      {stage037[27]},
      {stage037[171]}
   );
   gpc1_1 gpc1_1_1264(
      {stage037[28]},
      {stage037[172]}
   );
   gpc1_1 gpc1_1_1265(
      {stage037[29]},
      {stage037[173]}
   );
   gpc1_1 gpc1_1_1266(
      {stage037[30]},
      {stage037[174]}
   );
   gpc1_1 gpc1_1_1267(
      {stage037[31]},
      {stage037[175]}
   );
   gpc1_1 gpc1_1_1268(
      {stage037[32]},
      {stage037[176]}
   );
   gpc1_1 gpc1_1_1269(
      {stage037[33]},
      {stage037[177]}
   );
   gpc1_1 gpc1_1_1270(
      {stage037[34]},
      {stage037[178]}
   );
   gpc1_1 gpc1_1_1271(
      {stage037[35]},
      {stage037[179]}
   );
   gpc1_1 gpc1_1_1272(
      {stage037[36]},
      {stage037[180]}
   );
   gpc1_1 gpc1_1_1273(
      {stage037[37]},
      {stage037[181]}
   );
   gpc1_1 gpc1_1_1274(
      {stage037[38]},
      {stage037[182]}
   );
   gpc1_1 gpc1_1_1275(
      {stage037[39]},
      {stage037[183]}
   );
   gpc1_1 gpc1_1_1276(
      {stage037[40]},
      {stage037[184]}
   );
   gpc606_5 gpc606_5_1277(
      {stage037[41], stage037[42], stage037[43], stage037[44], stage037[45], stage037[46]},
      {stage039[0], stage039[1], stage039[2], stage039[3], stage039[4], stage039[5]},
      {stage041[128], stage040[138], stage039[141], stage038[151], stage037[185]}
   );
   gpc606_5 gpc606_5_1278(
      {stage037[47], stage037[48], stage037[49], stage037[50], stage037[51], stage037[52]},
      {stage039[6], stage039[7], stage039[8], stage039[9], stage039[10], stage039[11]},
      {stage041[129], stage040[139], stage039[142], stage038[152], stage037[186]}
   );
   gpc606_5 gpc606_5_1279(
      {stage037[53], stage037[54], stage037[55], stage037[56], stage037[57], stage037[58]},
      {stage039[12], stage039[13], stage039[14], stage039[15], stage039[16], stage039[17]},
      {stage041[130], stage040[140], stage039[143], stage038[153], stage037[187]}
   );
   gpc606_5 gpc606_5_1280(
      {stage037[59], stage037[60], stage037[61], stage037[62], stage037[63], stage037[64]},
      {stage039[18], stage039[19], stage039[20], stage039[21], stage039[22], stage039[23]},
      {stage041[131], stage040[141], stage039[144], stage038[154], stage037[188]}
   );
   gpc606_5 gpc606_5_1281(
      {stage037[65], stage037[66], stage037[67], stage037[68], stage037[69], stage037[70]},
      {stage039[24], stage039[25], stage039[26], stage039[27], stage039[28], stage039[29]},
      {stage041[132], stage040[142], stage039[145], stage038[155], stage037[189]}
   );
   gpc606_5 gpc606_5_1282(
      {stage037[71], stage037[72], stage037[73], stage037[74], stage037[75], stage037[76]},
      {stage039[30], stage039[31], stage039[32], stage039[33], stage039[34], stage039[35]},
      {stage041[133], stage040[143], stage039[146], stage038[156], stage037[190]}
   );
   gpc606_5 gpc606_5_1283(
      {stage037[77], stage037[78], stage037[79], stage037[80], stage037[81], stage037[82]},
      {stage039[36], stage039[37], stage039[38], stage039[39], stage039[40], stage039[41]},
      {stage041[134], stage040[144], stage039[147], stage038[157], stage037[191]}
   );
   gpc606_5 gpc606_5_1284(
      {stage037[83], stage037[84], stage037[85], stage037[86], stage037[87], stage037[88]},
      {stage039[42], stage039[43], stage039[44], stage039[45], stage039[46], stage039[47]},
      {stage041[135], stage040[145], stage039[148], stage038[158], stage037[192]}
   );
   gpc606_5 gpc606_5_1285(
      {stage037[89], stage037[90], stage037[91], stage037[92], stage037[93], stage037[94]},
      {stage039[48], stage039[49], stage039[50], stage039[51], stage039[52], stage039[53]},
      {stage041[136], stage040[146], stage039[149], stage038[159], stage037[193]}
   );
   gpc606_5 gpc606_5_1286(
      {stage037[95], stage037[96], stage037[97], stage037[98], stage037[99], stage037[100]},
      {stage039[54], stage039[55], stage039[56], stage039[57], stage039[58], stage039[59]},
      {stage041[137], stage040[147], stage039[150], stage038[160], stage037[194]}
   );
   gpc606_5 gpc606_5_1287(
      {stage037[101], stage037[102], stage037[103], stage037[104], stage037[105], stage037[106]},
      {stage039[60], stage039[61], stage039[62], stage039[63], stage039[64], stage039[65]},
      {stage041[138], stage040[148], stage039[151], stage038[161], stage037[195]}
   );
   gpc606_5 gpc606_5_1288(
      {stage037[107], stage037[108], stage037[109], stage037[110], stage037[111], stage037[112]},
      {stage039[66], stage039[67], stage039[68], stage039[69], stage039[70], stage039[71]},
      {stage041[139], stage040[149], stage039[152], stage038[162], stage037[196]}
   );
   gpc615_5 gpc615_5_1289(
      {stage037[113], stage037[114], stage037[115], stage037[116], stage037[117]},
      {stage038[62]},
      {stage039[72], stage039[73], stage039[74], stage039[75], stage039[76], stage039[77]},
      {stage041[140], stage040[150], stage039[153], stage038[163], stage037[197]}
   );
   gpc615_5 gpc615_5_1290(
      {stage037[118], stage037[119], stage037[120], stage037[121], stage037[122]},
      {stage038[63]},
      {stage039[78], stage039[79], stage039[80], stage039[81], stage039[82], stage039[83]},
      {stage041[141], stage040[151], stage039[154], stage038[164], stage037[198]}
   );
   gpc615_5 gpc615_5_1291(
      {stage037[123], stage037[124], stage037[125], stage037[126], stage037[127]},
      {stage038[64]},
      {stage039[84], stage039[85], stage039[86], stage039[87], stage039[88], stage039[89]},
      {stage041[142], stage040[152], stage039[155], stage038[165], stage037[199]}
   );
   gpc1_1 gpc1_1_1292(
      {stage038[65]},
      {stage038[166]}
   );
   gpc1_1 gpc1_1_1293(
      {stage038[66]},
      {stage038[167]}
   );
   gpc1_1 gpc1_1_1294(
      {stage038[67]},
      {stage038[168]}
   );
   gpc1_1 gpc1_1_1295(
      {stage038[68]},
      {stage038[169]}
   );
   gpc1_1 gpc1_1_1296(
      {stage038[69]},
      {stage038[170]}
   );
   gpc1_1 gpc1_1_1297(
      {stage038[70]},
      {stage038[171]}
   );
   gpc1_1 gpc1_1_1298(
      {stage038[71]},
      {stage038[172]}
   );
   gpc1_1 gpc1_1_1299(
      {stage038[72]},
      {stage038[173]}
   );
   gpc1_1 gpc1_1_1300(
      {stage038[73]},
      {stage038[174]}
   );
   gpc1_1 gpc1_1_1301(
      {stage038[74]},
      {stage038[175]}
   );
   gpc1_1 gpc1_1_1302(
      {stage038[75]},
      {stage038[176]}
   );
   gpc1_1 gpc1_1_1303(
      {stage038[76]},
      {stage038[177]}
   );
   gpc1_1 gpc1_1_1304(
      {stage038[77]},
      {stage038[178]}
   );
   gpc1_1 gpc1_1_1305(
      {stage038[78]},
      {stage038[179]}
   );
   gpc1_1 gpc1_1_1306(
      {stage038[79]},
      {stage038[180]}
   );
   gpc1_1 gpc1_1_1307(
      {stage038[80]},
      {stage038[181]}
   );
   gpc1_1 gpc1_1_1308(
      {stage038[81]},
      {stage038[182]}
   );
   gpc1_1 gpc1_1_1309(
      {stage038[82]},
      {stage038[183]}
   );
   gpc615_5 gpc615_5_1310(
      {stage038[83], stage038[84], stage038[85], stage038[86], stage038[87]},
      {stage039[90]},
      {stage040[0], stage040[1], stage040[2], stage040[3], stage040[4], stage040[5]},
      {stage042[128], stage041[143], stage040[153], stage039[156], stage038[184]}
   );
   gpc615_5 gpc615_5_1311(
      {stage038[88], stage038[89], stage038[90], stage038[91], stage038[92]},
      {stage039[91]},
      {stage040[6], stage040[7], stage040[8], stage040[9], stage040[10], stage040[11]},
      {stage042[129], stage041[144], stage040[154], stage039[157], stage038[185]}
   );
   gpc615_5 gpc615_5_1312(
      {stage038[93], stage038[94], stage038[95], stage038[96], stage038[97]},
      {stage039[92]},
      {stage040[12], stage040[13], stage040[14], stage040[15], stage040[16], stage040[17]},
      {stage042[130], stage041[145], stage040[155], stage039[158], stage038[186]}
   );
   gpc615_5 gpc615_5_1313(
      {stage038[98], stage038[99], stage038[100], stage038[101], stage038[102]},
      {stage039[93]},
      {stage040[18], stage040[19], stage040[20], stage040[21], stage040[22], stage040[23]},
      {stage042[131], stage041[146], stage040[156], stage039[159], stage038[187]}
   );
   gpc615_5 gpc615_5_1314(
      {stage038[103], stage038[104], stage038[105], stage038[106], stage038[107]},
      {stage039[94]},
      {stage040[24], stage040[25], stage040[26], stage040[27], stage040[28], stage040[29]},
      {stage042[132], stage041[147], stage040[157], stage039[160], stage038[188]}
   );
   gpc615_5 gpc615_5_1315(
      {stage038[108], stage038[109], stage038[110], stage038[111], stage038[112]},
      {stage039[95]},
      {stage040[30], stage040[31], stage040[32], stage040[33], stage040[34], stage040[35]},
      {stage042[133], stage041[148], stage040[158], stage039[161], stage038[189]}
   );
   gpc615_5 gpc615_5_1316(
      {stage038[113], stage038[114], stage038[115], stage038[116], stage038[117]},
      {stage039[96]},
      {stage040[36], stage040[37], stage040[38], stage040[39], stage040[40], stage040[41]},
      {stage042[134], stage041[149], stage040[159], stage039[162], stage038[190]}
   );
   gpc615_5 gpc615_5_1317(
      {stage038[118], stage038[119], stage038[120], stage038[121], stage038[122]},
      {stage039[97]},
      {stage040[42], stage040[43], stage040[44], stage040[45], stage040[46], stage040[47]},
      {stage042[135], stage041[150], stage040[160], stage039[163], stage038[191]}
   );
   gpc615_5 gpc615_5_1318(
      {stage038[123], stage038[124], stage038[125], stage038[126], stage038[127]},
      {stage039[98]},
      {stage040[48], stage040[49], stage040[50], stage040[51], stage040[52], stage040[53]},
      {stage042[136], stage041[151], stage040[161], stage039[164], stage038[192]}
   );
   gpc1_1 gpc1_1_1319(
      {stage039[99]},
      {stage039[165]}
   );
   gpc1_1 gpc1_1_1320(
      {stage039[100]},
      {stage039[166]}
   );
   gpc1_1 gpc1_1_1321(
      {stage039[101]},
      {stage039[167]}
   );
   gpc1_1 gpc1_1_1322(
      {stage039[102]},
      {stage039[168]}
   );
   gpc1_1 gpc1_1_1323(
      {stage039[103]},
      {stage039[169]}
   );
   gpc1_1 gpc1_1_1324(
      {stage039[104]},
      {stage039[170]}
   );
   gpc1_1 gpc1_1_1325(
      {stage039[105]},
      {stage039[171]}
   );
   gpc1_1 gpc1_1_1326(
      {stage039[106]},
      {stage039[172]}
   );
   gpc1_1 gpc1_1_1327(
      {stage039[107]},
      {stage039[173]}
   );
   gpc1_1 gpc1_1_1328(
      {stage039[108]},
      {stage039[174]}
   );
   gpc1_1 gpc1_1_1329(
      {stage039[109]},
      {stage039[175]}
   );
   gpc1_1 gpc1_1_1330(
      {stage039[110]},
      {stage039[176]}
   );
   gpc1_1 gpc1_1_1331(
      {stage039[111]},
      {stage039[177]}
   );
   gpc1_1 gpc1_1_1332(
      {stage039[112]},
      {stage039[178]}
   );
   gpc1_1 gpc1_1_1333(
      {stage039[113]},
      {stage039[179]}
   );
   gpc1_1 gpc1_1_1334(
      {stage039[114]},
      {stage039[180]}
   );
   gpc1_1 gpc1_1_1335(
      {stage039[115]},
      {stage039[181]}
   );
   gpc1_1 gpc1_1_1336(
      {stage039[116]},
      {stage039[182]}
   );
   gpc1_1 gpc1_1_1337(
      {stage039[117]},
      {stage039[183]}
   );
   gpc1_1 gpc1_1_1338(
      {stage039[118]},
      {stage039[184]}
   );
   gpc1_1 gpc1_1_1339(
      {stage039[119]},
      {stage039[185]}
   );
   gpc1_1 gpc1_1_1340(
      {stage039[120]},
      {stage039[186]}
   );
   gpc1_1 gpc1_1_1341(
      {stage039[121]},
      {stage039[187]}
   );
   gpc606_5 gpc606_5_1342(
      {stage039[122], stage039[123], stage039[124], stage039[125], stage039[126], stage039[127]},
      {stage041[0], stage041[1], stage041[2], stage041[3], stage041[4], stage041[5]},
      {stage043[128], stage042[137], stage041[152], stage040[162], stage039[188]}
   );
   gpc1_1 gpc1_1_1343(
      {stage040[54]},
      {stage040[163]}
   );
   gpc1_1 gpc1_1_1344(
      {stage040[55]},
      {stage040[164]}
   );
   gpc1_1 gpc1_1_1345(
      {stage040[56]},
      {stage040[165]}
   );
   gpc1_1 gpc1_1_1346(
      {stage040[57]},
      {stage040[166]}
   );
   gpc1_1 gpc1_1_1347(
      {stage040[58]},
      {stage040[167]}
   );
   gpc1_1 gpc1_1_1348(
      {stage040[59]},
      {stage040[168]}
   );
   gpc1_1 gpc1_1_1349(
      {stage040[60]},
      {stage040[169]}
   );
   gpc1_1 gpc1_1_1350(
      {stage040[61]},
      {stage040[170]}
   );
   gpc1_1 gpc1_1_1351(
      {stage040[62]},
      {stage040[171]}
   );
   gpc1_1 gpc1_1_1352(
      {stage040[63]},
      {stage040[172]}
   );
   gpc1_1 gpc1_1_1353(
      {stage040[64]},
      {stage040[173]}
   );
   gpc1_1 gpc1_1_1354(
      {stage040[65]},
      {stage040[174]}
   );
   gpc1_1 gpc1_1_1355(
      {stage040[66]},
      {stage040[175]}
   );
   gpc1_1 gpc1_1_1356(
      {stage040[67]},
      {stage040[176]}
   );
   gpc1_1 gpc1_1_1357(
      {stage040[68]},
      {stage040[177]}
   );
   gpc1_1 gpc1_1_1358(
      {stage040[69]},
      {stage040[178]}
   );
   gpc1_1 gpc1_1_1359(
      {stage040[70]},
      {stage040[179]}
   );
   gpc1_1 gpc1_1_1360(
      {stage040[71]},
      {stage040[180]}
   );
   gpc1_1 gpc1_1_1361(
      {stage040[72]},
      {stage040[181]}
   );
   gpc1_1 gpc1_1_1362(
      {stage040[73]},
      {stage040[182]}
   );
   gpc1_1 gpc1_1_1363(
      {stage040[74]},
      {stage040[183]}
   );
   gpc1_1 gpc1_1_1364(
      {stage040[75]},
      {stage040[184]}
   );
   gpc1_1 gpc1_1_1365(
      {stage040[76]},
      {stage040[185]}
   );
   gpc1_1 gpc1_1_1366(
      {stage040[77]},
      {stage040[186]}
   );
   gpc1_1 gpc1_1_1367(
      {stage040[78]},
      {stage040[187]}
   );
   gpc1_1 gpc1_1_1368(
      {stage040[79]},
      {stage040[188]}
   );
   gpc1_1 gpc1_1_1369(
      {stage040[80]},
      {stage040[189]}
   );
   gpc1_1 gpc1_1_1370(
      {stage040[81]},
      {stage040[190]}
   );
   gpc1_1 gpc1_1_1371(
      {stage040[82]},
      {stage040[191]}
   );
   gpc1_1 gpc1_1_1372(
      {stage040[83]},
      {stage040[192]}
   );
   gpc1_1 gpc1_1_1373(
      {stage040[84]},
      {stage040[193]}
   );
   gpc1_1 gpc1_1_1374(
      {stage040[85]},
      {stage040[194]}
   );
   gpc1_1 gpc1_1_1375(
      {stage040[86]},
      {stage040[195]}
   );
   gpc1_1 gpc1_1_1376(
      {stage040[87]},
      {stage040[196]}
   );
   gpc1_1 gpc1_1_1377(
      {stage040[88]},
      {stage040[197]}
   );
   gpc1_1 gpc1_1_1378(
      {stage040[89]},
      {stage040[198]}
   );
   gpc1_1 gpc1_1_1379(
      {stage040[90]},
      {stage040[199]}
   );
   gpc1_1 gpc1_1_1380(
      {stage040[91]},
      {stage040[200]}
   );
   gpc1_1 gpc1_1_1381(
      {stage040[92]},
      {stage040[201]}
   );
   gpc1_1 gpc1_1_1382(
      {stage040[93]},
      {stage040[202]}
   );
   gpc1_1 gpc1_1_1383(
      {stage040[94]},
      {stage040[203]}
   );
   gpc1_1 gpc1_1_1384(
      {stage040[95]},
      {stage040[204]}
   );
   gpc1_1 gpc1_1_1385(
      {stage040[96]},
      {stage040[205]}
   );
   gpc1_1 gpc1_1_1386(
      {stage040[97]},
      {stage040[206]}
   );
   gpc1_1 gpc1_1_1387(
      {stage040[98]},
      {stage040[207]}
   );
   gpc1_1 gpc1_1_1388(
      {stage040[99]},
      {stage040[208]}
   );
   gpc1_1 gpc1_1_1389(
      {stage040[100]},
      {stage040[209]}
   );
   gpc1_1 gpc1_1_1390(
      {stage040[101]},
      {stage040[210]}
   );
   gpc1_1 gpc1_1_1391(
      {stage040[102]},
      {stage040[211]}
   );
   gpc1_1 gpc1_1_1392(
      {stage040[103]},
      {stage040[212]}
   );
   gpc1_1 gpc1_1_1393(
      {stage040[104]},
      {stage040[213]}
   );
   gpc606_5 gpc606_5_1394(
      {stage040[105], stage040[106], stage040[107], stage040[108], stage040[109], stage040[110]},
      {stage042[0], stage042[1], stage042[2], stage042[3], stage042[4], stage042[5]},
      {stage044[128], stage043[129], stage042[138], stage041[153], stage040[214]}
   );
   gpc606_5 gpc606_5_1395(
      {stage040[111], stage040[112], stage040[113], stage040[114], stage040[115], stage040[116]},
      {stage042[6], stage042[7], stage042[8], stage042[9], stage042[10], stage042[11]},
      {stage044[129], stage043[130], stage042[139], stage041[154], stage040[215]}
   );
   gpc606_5 gpc606_5_1396(
      {stage040[117], stage040[118], stage040[119], stage040[120], stage040[121], stage040[122]},
      {stage042[12], stage042[13], stage042[14], stage042[15], stage042[16], stage042[17]},
      {stage044[130], stage043[131], stage042[140], stage041[155], stage040[216]}
   );
   gpc2135_5 gpc2135_5_1397(
      {stage040[123], stage040[124], stage040[125], stage040[126], stage040[127]},
      {stage041[6], stage041[7], stage041[8]},
      {stage042[18]},
      {stage043[0], stage043[1]},
      {stage044[131], stage043[132], stage042[141], stage041[156], stage040[217]}
   );
   gpc1_1 gpc1_1_1398(
      {stage041[9]},
      {stage041[157]}
   );
   gpc1_1 gpc1_1_1399(
      {stage041[10]},
      {stage041[158]}
   );
   gpc1_1 gpc1_1_1400(
      {stage041[11]},
      {stage041[159]}
   );
   gpc1_1 gpc1_1_1401(
      {stage041[12]},
      {stage041[160]}
   );
   gpc1_1 gpc1_1_1402(
      {stage041[13]},
      {stage041[161]}
   );
   gpc1_1 gpc1_1_1403(
      {stage041[14]},
      {stage041[162]}
   );
   gpc1_1 gpc1_1_1404(
      {stage041[15]},
      {stage041[163]}
   );
   gpc1_1 gpc1_1_1405(
      {stage041[16]},
      {stage041[164]}
   );
   gpc1_1 gpc1_1_1406(
      {stage041[17]},
      {stage041[165]}
   );
   gpc1_1 gpc1_1_1407(
      {stage041[18]},
      {stage041[166]}
   );
   gpc1_1 gpc1_1_1408(
      {stage041[19]},
      {stage041[167]}
   );
   gpc1_1 gpc1_1_1409(
      {stage041[20]},
      {stage041[168]}
   );
   gpc1_1 gpc1_1_1410(
      {stage041[21]},
      {stage041[169]}
   );
   gpc1_1 gpc1_1_1411(
      {stage041[22]},
      {stage041[170]}
   );
   gpc1_1 gpc1_1_1412(
      {stage041[23]},
      {stage041[171]}
   );
   gpc1_1 gpc1_1_1413(
      {stage041[24]},
      {stage041[172]}
   );
   gpc1_1 gpc1_1_1414(
      {stage041[25]},
      {stage041[173]}
   );
   gpc1_1 gpc1_1_1415(
      {stage041[26]},
      {stage041[174]}
   );
   gpc1_1 gpc1_1_1416(
      {stage041[27]},
      {stage041[175]}
   );
   gpc1_1 gpc1_1_1417(
      {stage041[28]},
      {stage041[176]}
   );
   gpc1_1 gpc1_1_1418(
      {stage041[29]},
      {stage041[177]}
   );
   gpc1_1 gpc1_1_1419(
      {stage041[30]},
      {stage041[178]}
   );
   gpc1_1 gpc1_1_1420(
      {stage041[31]},
      {stage041[179]}
   );
   gpc1_1 gpc1_1_1421(
      {stage041[32]},
      {stage041[180]}
   );
   gpc1_1 gpc1_1_1422(
      {stage041[33]},
      {stage041[181]}
   );
   gpc1_1 gpc1_1_1423(
      {stage041[34]},
      {stage041[182]}
   );
   gpc1_1 gpc1_1_1424(
      {stage041[35]},
      {stage041[183]}
   );
   gpc1_1 gpc1_1_1425(
      {stage041[36]},
      {stage041[184]}
   );
   gpc606_5 gpc606_5_1426(
      {stage041[37], stage041[38], stage041[39], stage041[40], stage041[41], stage041[42]},
      {stage043[2], stage043[3], stage043[4], stage043[5], stage043[6], stage043[7]},
      {stage045[128], stage044[132], stage043[133], stage042[142], stage041[185]}
   );
   gpc606_5 gpc606_5_1427(
      {stage041[43], stage041[44], stage041[45], stage041[46], stage041[47], stage041[48]},
      {stage043[8], stage043[9], stage043[10], stage043[11], stage043[12], stage043[13]},
      {stage045[129], stage044[133], stage043[134], stage042[143], stage041[186]}
   );
   gpc606_5 gpc606_5_1428(
      {stage041[49], stage041[50], stage041[51], stage041[52], stage041[53], stage041[54]},
      {stage043[14], stage043[15], stage043[16], stage043[17], stage043[18], stage043[19]},
      {stage045[130], stage044[134], stage043[135], stage042[144], stage041[187]}
   );
   gpc606_5 gpc606_5_1429(
      {stage041[55], stage041[56], stage041[57], stage041[58], stage041[59], stage041[60]},
      {stage043[20], stage043[21], stage043[22], stage043[23], stage043[24], stage043[25]},
      {stage045[131], stage044[135], stage043[136], stage042[145], stage041[188]}
   );
   gpc606_5 gpc606_5_1430(
      {stage041[61], stage041[62], stage041[63], stage041[64], stage041[65], stage041[66]},
      {stage043[26], stage043[27], stage043[28], stage043[29], stage043[30], stage043[31]},
      {stage045[132], stage044[136], stage043[137], stage042[146], stage041[189]}
   );
   gpc606_5 gpc606_5_1431(
      {stage041[67], stage041[68], stage041[69], stage041[70], stage041[71], stage041[72]},
      {stage043[32], stage043[33], stage043[34], stage043[35], stage043[36], stage043[37]},
      {stage045[133], stage044[137], stage043[138], stage042[147], stage041[190]}
   );
   gpc615_5 gpc615_5_1432(
      {stage041[73], stage041[74], stage041[75], stage041[76], stage041[77]},
      {stage042[19]},
      {stage043[38], stage043[39], stage043[40], stage043[41], stage043[42], stage043[43]},
      {stage045[134], stage044[138], stage043[139], stage042[148], stage041[191]}
   );
   gpc615_5 gpc615_5_1433(
      {stage041[78], stage041[79], stage041[80], stage041[81], stage041[82]},
      {stage042[20]},
      {stage043[44], stage043[45], stage043[46], stage043[47], stage043[48], stage043[49]},
      {stage045[135], stage044[139], stage043[140], stage042[149], stage041[192]}
   );
   gpc615_5 gpc615_5_1434(
      {stage041[83], stage041[84], stage041[85], stage041[86], stage041[87]},
      {stage042[21]},
      {stage043[50], stage043[51], stage043[52], stage043[53], stage043[54], stage043[55]},
      {stage045[136], stage044[140], stage043[141], stage042[150], stage041[193]}
   );
   gpc615_5 gpc615_5_1435(
      {stage041[88], stage041[89], stage041[90], stage041[91], stage041[92]},
      {stage042[22]},
      {stage043[56], stage043[57], stage043[58], stage043[59], stage043[60], stage043[61]},
      {stage045[137], stage044[141], stage043[142], stage042[151], stage041[194]}
   );
   gpc615_5 gpc615_5_1436(
      {stage041[93], stage041[94], stage041[95], stage041[96], stage041[97]},
      {stage042[23]},
      {stage043[62], stage043[63], stage043[64], stage043[65], stage043[66], stage043[67]},
      {stage045[138], stage044[142], stage043[143], stage042[152], stage041[195]}
   );
   gpc615_5 gpc615_5_1437(
      {stage041[98], stage041[99], stage041[100], stage041[101], stage041[102]},
      {stage042[24]},
      {stage043[68], stage043[69], stage043[70], stage043[71], stage043[72], stage043[73]},
      {stage045[139], stage044[143], stage043[144], stage042[153], stage041[196]}
   );
   gpc615_5 gpc615_5_1438(
      {stage041[103], stage041[104], stage041[105], stage041[106], stage041[107]},
      {stage042[25]},
      {stage043[74], stage043[75], stage043[76], stage043[77], stage043[78], stage043[79]},
      {stage045[140], stage044[144], stage043[145], stage042[154], stage041[197]}
   );
   gpc615_5 gpc615_5_1439(
      {stage041[108], stage041[109], stage041[110], stage041[111], stage041[112]},
      {stage042[26]},
      {stage043[80], stage043[81], stage043[82], stage043[83], stage043[84], stage043[85]},
      {stage045[141], stage044[145], stage043[146], stage042[155], stage041[198]}
   );
   gpc615_5 gpc615_5_1440(
      {stage041[113], stage041[114], stage041[115], stage041[116], stage041[117]},
      {stage042[27]},
      {stage043[86], stage043[87], stage043[88], stage043[89], stage043[90], stage043[91]},
      {stage045[142], stage044[146], stage043[147], stage042[156], stage041[199]}
   );
   gpc615_5 gpc615_5_1441(
      {stage041[118], stage041[119], stage041[120], stage041[121], stage041[122]},
      {stage042[28]},
      {stage043[92], stage043[93], stage043[94], stage043[95], stage043[96], stage043[97]},
      {stage045[143], stage044[147], stage043[148], stage042[157], stage041[200]}
   );
   gpc615_5 gpc615_5_1442(
      {stage041[123], stage041[124], stage041[125], stage041[126], stage041[127]},
      {stage042[29]},
      {stage043[98], stage043[99], stage043[100], stage043[101], stage043[102], stage043[103]},
      {stage045[144], stage044[148], stage043[149], stage042[158], stage041[201]}
   );
   gpc1_1 gpc1_1_1443(
      {stage042[30]},
      {stage042[159]}
   );
   gpc1_1 gpc1_1_1444(
      {stage042[31]},
      {stage042[160]}
   );
   gpc1_1 gpc1_1_1445(
      {stage042[32]},
      {stage042[161]}
   );
   gpc1_1 gpc1_1_1446(
      {stage042[33]},
      {stage042[162]}
   );
   gpc1_1 gpc1_1_1447(
      {stage042[34]},
      {stage042[163]}
   );
   gpc1_1 gpc1_1_1448(
      {stage042[35]},
      {stage042[164]}
   );
   gpc1_1 gpc1_1_1449(
      {stage042[36]},
      {stage042[165]}
   );
   gpc1_1 gpc1_1_1450(
      {stage042[37]},
      {stage042[166]}
   );
   gpc1_1 gpc1_1_1451(
      {stage042[38]},
      {stage042[167]}
   );
   gpc1_1 gpc1_1_1452(
      {stage042[39]},
      {stage042[168]}
   );
   gpc1_1 gpc1_1_1453(
      {stage042[40]},
      {stage042[169]}
   );
   gpc1_1 gpc1_1_1454(
      {stage042[41]},
      {stage042[170]}
   );
   gpc1_1 gpc1_1_1455(
      {stage042[42]},
      {stage042[171]}
   );
   gpc1_1 gpc1_1_1456(
      {stage042[43]},
      {stage042[172]}
   );
   gpc1_1 gpc1_1_1457(
      {stage042[44]},
      {stage042[173]}
   );
   gpc1_1 gpc1_1_1458(
      {stage042[45]},
      {stage042[174]}
   );
   gpc1_1 gpc1_1_1459(
      {stage042[46]},
      {stage042[175]}
   );
   gpc1_1 gpc1_1_1460(
      {stage042[47]},
      {stage042[176]}
   );
   gpc1_1 gpc1_1_1461(
      {stage042[48]},
      {stage042[177]}
   );
   gpc1_1 gpc1_1_1462(
      {stage042[49]},
      {stage042[178]}
   );
   gpc1_1 gpc1_1_1463(
      {stage042[50]},
      {stage042[179]}
   );
   gpc1_1 gpc1_1_1464(
      {stage042[51]},
      {stage042[180]}
   );
   gpc1_1 gpc1_1_1465(
      {stage042[52]},
      {stage042[181]}
   );
   gpc1_1 gpc1_1_1466(
      {stage042[53]},
      {stage042[182]}
   );
   gpc1_1 gpc1_1_1467(
      {stage042[54]},
      {stage042[183]}
   );
   gpc1_1 gpc1_1_1468(
      {stage042[55]},
      {stage042[184]}
   );
   gpc1_1 gpc1_1_1469(
      {stage042[56]},
      {stage042[185]}
   );
   gpc1_1 gpc1_1_1470(
      {stage042[57]},
      {stage042[186]}
   );
   gpc1_1 gpc1_1_1471(
      {stage042[58]},
      {stage042[187]}
   );
   gpc1_1 gpc1_1_1472(
      {stage042[59]},
      {stage042[188]}
   );
   gpc1_1 gpc1_1_1473(
      {stage042[60]},
      {stage042[189]}
   );
   gpc1_1 gpc1_1_1474(
      {stage042[61]},
      {stage042[190]}
   );
   gpc1_1 gpc1_1_1475(
      {stage042[62]},
      {stage042[191]}
   );
   gpc1_1 gpc1_1_1476(
      {stage042[63]},
      {stage042[192]}
   );
   gpc1_1 gpc1_1_1477(
      {stage042[64]},
      {stage042[193]}
   );
   gpc1_1 gpc1_1_1478(
      {stage042[65]},
      {stage042[194]}
   );
   gpc1_1 gpc1_1_1479(
      {stage042[66]},
      {stage042[195]}
   );
   gpc1_1 gpc1_1_1480(
      {stage042[67]},
      {stage042[196]}
   );
   gpc615_5 gpc615_5_1481(
      {stage042[68], stage042[69], stage042[70], stage042[71], stage042[72]},
      {stage043[104]},
      {stage044[0], stage044[1], stage044[2], stage044[3], stage044[4], stage044[5]},
      {stage046[128], stage045[145], stage044[149], stage043[150], stage042[197]}
   );
   gpc615_5 gpc615_5_1482(
      {stage042[73], stage042[74], stage042[75], stage042[76], stage042[77]},
      {stage043[105]},
      {stage044[6], stage044[7], stage044[8], stage044[9], stage044[10], stage044[11]},
      {stage046[129], stage045[146], stage044[150], stage043[151], stage042[198]}
   );
   gpc615_5 gpc615_5_1483(
      {stage042[78], stage042[79], stage042[80], stage042[81], stage042[82]},
      {stage043[106]},
      {stage044[12], stage044[13], stage044[14], stage044[15], stage044[16], stage044[17]},
      {stage046[130], stage045[147], stage044[151], stage043[152], stage042[199]}
   );
   gpc615_5 gpc615_5_1484(
      {stage042[83], stage042[84], stage042[85], stage042[86], stage042[87]},
      {stage043[107]},
      {stage044[18], stage044[19], stage044[20], stage044[21], stage044[22], stage044[23]},
      {stage046[131], stage045[148], stage044[152], stage043[153], stage042[200]}
   );
   gpc615_5 gpc615_5_1485(
      {stage042[88], stage042[89], stage042[90], stage042[91], stage042[92]},
      {stage043[108]},
      {stage044[24], stage044[25], stage044[26], stage044[27], stage044[28], stage044[29]},
      {stage046[132], stage045[149], stage044[153], stage043[154], stage042[201]}
   );
   gpc615_5 gpc615_5_1486(
      {stage042[93], stage042[94], stage042[95], stage042[96], stage042[97]},
      {stage043[109]},
      {stage044[30], stage044[31], stage044[32], stage044[33], stage044[34], stage044[35]},
      {stage046[133], stage045[150], stage044[154], stage043[155], stage042[202]}
   );
   gpc615_5 gpc615_5_1487(
      {stage042[98], stage042[99], stage042[100], stage042[101], stage042[102]},
      {stage043[110]},
      {stage044[36], stage044[37], stage044[38], stage044[39], stage044[40], stage044[41]},
      {stage046[134], stage045[151], stage044[155], stage043[156], stage042[203]}
   );
   gpc615_5 gpc615_5_1488(
      {stage042[103], stage042[104], stage042[105], stage042[106], stage042[107]},
      {stage043[111]},
      {stage044[42], stage044[43], stage044[44], stage044[45], stage044[46], stage044[47]},
      {stage046[135], stage045[152], stage044[156], stage043[157], stage042[204]}
   );
   gpc615_5 gpc615_5_1489(
      {stage042[108], stage042[109], stage042[110], stage042[111], stage042[112]},
      {stage043[112]},
      {stage044[48], stage044[49], stage044[50], stage044[51], stage044[52], stage044[53]},
      {stage046[136], stage045[153], stage044[157], stage043[158], stage042[205]}
   );
   gpc615_5 gpc615_5_1490(
      {stage042[113], stage042[114], stage042[115], stage042[116], stage042[117]},
      {stage043[113]},
      {stage044[54], stage044[55], stage044[56], stage044[57], stage044[58], stage044[59]},
      {stage046[137], stage045[154], stage044[158], stage043[159], stage042[206]}
   );
   gpc615_5 gpc615_5_1491(
      {stage042[118], stage042[119], stage042[120], stage042[121], stage042[122]},
      {stage043[114]},
      {stage044[60], stage044[61], stage044[62], stage044[63], stage044[64], stage044[65]},
      {stage046[138], stage045[155], stage044[159], stage043[160], stage042[207]}
   );
   gpc615_5 gpc615_5_1492(
      {stage042[123], stage042[124], stage042[125], stage042[126], stage042[127]},
      {stage043[115]},
      {stage044[66], stage044[67], stage044[68], stage044[69], stage044[70], stage044[71]},
      {stage046[139], stage045[156], stage044[160], stage043[161], stage042[208]}
   );
   gpc1_1 gpc1_1_1493(
      {stage043[116]},
      {stage043[162]}
   );
   gpc1_1 gpc1_1_1494(
      {stage043[117]},
      {stage043[163]}
   );
   gpc615_5 gpc615_5_1495(
      {stage043[118], stage043[119], stage043[120], stage043[121], stage043[122]},
      {stage044[72]},
      {stage045[0], stage045[1], stage045[2], stage045[3], stage045[4], stage045[5]},
      {stage047[128], stage046[140], stage045[157], stage044[161], stage043[164]}
   );
   gpc615_5 gpc615_5_1496(
      {stage043[123], stage043[124], stage043[125], stage043[126], stage043[127]},
      {stage044[73]},
      {stage045[6], stage045[7], stage045[8], stage045[9], stage045[10], stage045[11]},
      {stage047[129], stage046[141], stage045[158], stage044[162], stage043[165]}
   );
   gpc1_1 gpc1_1_1497(
      {stage044[74]},
      {stage044[163]}
   );
   gpc1_1 gpc1_1_1498(
      {stage044[75]},
      {stage044[164]}
   );
   gpc1_1 gpc1_1_1499(
      {stage044[76]},
      {stage044[165]}
   );
   gpc1_1 gpc1_1_1500(
      {stage044[77]},
      {stage044[166]}
   );
   gpc1_1 gpc1_1_1501(
      {stage044[78]},
      {stage044[167]}
   );
   gpc1_1 gpc1_1_1502(
      {stage044[79]},
      {stage044[168]}
   );
   gpc1_1 gpc1_1_1503(
      {stage044[80]},
      {stage044[169]}
   );
   gpc1_1 gpc1_1_1504(
      {stage044[81]},
      {stage044[170]}
   );
   gpc606_5 gpc606_5_1505(
      {stage044[82], stage044[83], stage044[84], stage044[85], stage044[86], stage044[87]},
      {stage046[0], stage046[1], stage046[2], stage046[3], stage046[4], stage046[5]},
      {stage048[128], stage047[130], stage046[142], stage045[159], stage044[171]}
   );
   gpc606_5 gpc606_5_1506(
      {stage044[88], stage044[89], stage044[90], stage044[91], stage044[92], stage044[93]},
      {stage046[6], stage046[7], stage046[8], stage046[9], stage046[10], stage046[11]},
      {stage048[129], stage047[131], stage046[143], stage045[160], stage044[172]}
   );
   gpc606_5 gpc606_5_1507(
      {stage044[94], stage044[95], stage044[96], stage044[97], stage044[98], stage044[99]},
      {stage046[12], stage046[13], stage046[14], stage046[15], stage046[16], stage046[17]},
      {stage048[130], stage047[132], stage046[144], stage045[161], stage044[173]}
   );
   gpc606_5 gpc606_5_1508(
      {stage044[100], stage044[101], stage044[102], stage044[103], stage044[104], stage044[105]},
      {stage046[18], stage046[19], stage046[20], stage046[21], stage046[22], stage046[23]},
      {stage048[131], stage047[133], stage046[145], stage045[162], stage044[174]}
   );
   gpc606_5 gpc606_5_1509(
      {stage044[106], stage044[107], stage044[108], stage044[109], stage044[110], stage044[111]},
      {stage046[24], stage046[25], stage046[26], stage046[27], stage046[28], stage046[29]},
      {stage048[132], stage047[134], stage046[146], stage045[163], stage044[175]}
   );
   gpc606_5 gpc606_5_1510(
      {stage044[112], stage044[113], stage044[114], stage044[115], stage044[116], stage044[117]},
      {stage046[30], stage046[31], stage046[32], stage046[33], stage046[34], stage046[35]},
      {stage048[133], stage047[135], stage046[147], stage045[164], stage044[176]}
   );
   gpc615_5 gpc615_5_1511(
      {stage044[118], stage044[119], stage044[120], stage044[121], stage044[122]},
      {stage045[12]},
      {stage046[36], stage046[37], stage046[38], stage046[39], stage046[40], stage046[41]},
      {stage048[134], stage047[136], stage046[148], stage045[165], stage044[177]}
   );
   gpc615_5 gpc615_5_1512(
      {stage044[123], stage044[124], stage044[125], stage044[126], stage044[127]},
      {stage045[13]},
      {stage046[42], stage046[43], stage046[44], stage046[45], stage046[46], stage046[47]},
      {stage048[135], stage047[137], stage046[149], stage045[166], stage044[178]}
   );
   gpc1_1 gpc1_1_1513(
      {stage045[14]},
      {stage045[167]}
   );
   gpc1_1 gpc1_1_1514(
      {stage045[15]},
      {stage045[168]}
   );
   gpc1_1 gpc1_1_1515(
      {stage045[16]},
      {stage045[169]}
   );
   gpc1_1 gpc1_1_1516(
      {stage045[17]},
      {stage045[170]}
   );
   gpc1_1 gpc1_1_1517(
      {stage045[18]},
      {stage045[171]}
   );
   gpc1_1 gpc1_1_1518(
      {stage045[19]},
      {stage045[172]}
   );
   gpc1_1 gpc1_1_1519(
      {stage045[20]},
      {stage045[173]}
   );
   gpc1_1 gpc1_1_1520(
      {stage045[21]},
      {stage045[174]}
   );
   gpc1_1 gpc1_1_1521(
      {stage045[22]},
      {stage045[175]}
   );
   gpc1_1 gpc1_1_1522(
      {stage045[23]},
      {stage045[176]}
   );
   gpc1_1 gpc1_1_1523(
      {stage045[24]},
      {stage045[177]}
   );
   gpc1_1 gpc1_1_1524(
      {stage045[25]},
      {stage045[178]}
   );
   gpc1_1 gpc1_1_1525(
      {stage045[26]},
      {stage045[179]}
   );
   gpc1_1 gpc1_1_1526(
      {stage045[27]},
      {stage045[180]}
   );
   gpc1_1 gpc1_1_1527(
      {stage045[28]},
      {stage045[181]}
   );
   gpc1_1 gpc1_1_1528(
      {stage045[29]},
      {stage045[182]}
   );
   gpc1_1 gpc1_1_1529(
      {stage045[30]},
      {stage045[183]}
   );
   gpc1_1 gpc1_1_1530(
      {stage045[31]},
      {stage045[184]}
   );
   gpc1_1 gpc1_1_1531(
      {stage045[32]},
      {stage045[185]}
   );
   gpc1_1 gpc1_1_1532(
      {stage045[33]},
      {stage045[186]}
   );
   gpc1_1 gpc1_1_1533(
      {stage045[34]},
      {stage045[187]}
   );
   gpc623_5 gpc623_5_1534(
      {stage045[35], stage045[36], stage045[37]},
      {stage046[48], stage046[49]},
      {stage047[0], stage047[1], stage047[2], stage047[3], stage047[4], stage047[5]},
      {stage049[128], stage048[136], stage047[138], stage046[150], stage045[188]}
   );
   gpc606_5 gpc606_5_1535(
      {stage045[38], stage045[39], stage045[40], stage045[41], stage045[42], stage045[43]},
      {stage047[6], stage047[7], stage047[8], stage047[9], stage047[10], stage047[11]},
      {stage049[129], stage048[137], stage047[139], stage046[151], stage045[189]}
   );
   gpc606_5 gpc606_5_1536(
      {stage045[44], stage045[45], stage045[46], stage045[47], stage045[48], stage045[49]},
      {stage047[12], stage047[13], stage047[14], stage047[15], stage047[16], stage047[17]},
      {stage049[130], stage048[138], stage047[140], stage046[152], stage045[190]}
   );
   gpc606_5 gpc606_5_1537(
      {stage045[50], stage045[51], stage045[52], stage045[53], stage045[54], stage045[55]},
      {stage047[18], stage047[19], stage047[20], stage047[21], stage047[22], stage047[23]},
      {stage049[131], stage048[139], stage047[141], stage046[153], stage045[191]}
   );
   gpc606_5 gpc606_5_1538(
      {stage045[56], stage045[57], stage045[58], stage045[59], stage045[60], stage045[61]},
      {stage047[24], stage047[25], stage047[26], stage047[27], stage047[28], stage047[29]},
      {stage049[132], stage048[140], stage047[142], stage046[154], stage045[192]}
   );
   gpc606_5 gpc606_5_1539(
      {stage045[62], stage045[63], stage045[64], stage045[65], stage045[66], stage045[67]},
      {stage047[30], stage047[31], stage047[32], stage047[33], stage047[34], stage047[35]},
      {stage049[133], stage048[141], stage047[143], stage046[155], stage045[193]}
   );
   gpc606_5 gpc606_5_1540(
      {stage045[68], stage045[69], stage045[70], stage045[71], stage045[72], stage045[73]},
      {stage047[36], stage047[37], stage047[38], stage047[39], stage047[40], stage047[41]},
      {stage049[134], stage048[142], stage047[144], stage046[156], stage045[194]}
   );
   gpc606_5 gpc606_5_1541(
      {stage045[74], stage045[75], stage045[76], stage045[77], stage045[78], stage045[79]},
      {stage047[42], stage047[43], stage047[44], stage047[45], stage047[46], stage047[47]},
      {stage049[135], stage048[143], stage047[145], stage046[157], stage045[195]}
   );
   gpc606_5 gpc606_5_1542(
      {stage045[80], stage045[81], stage045[82], stage045[83], stage045[84], stage045[85]},
      {stage047[48], stage047[49], stage047[50], stage047[51], stage047[52], stage047[53]},
      {stage049[136], stage048[144], stage047[146], stage046[158], stage045[196]}
   );
   gpc606_5 gpc606_5_1543(
      {stage045[86], stage045[87], stage045[88], stage045[89], stage045[90], stage045[91]},
      {stage047[54], stage047[55], stage047[56], stage047[57], stage047[58], stage047[59]},
      {stage049[137], stage048[145], stage047[147], stage046[159], stage045[197]}
   );
   gpc606_5 gpc606_5_1544(
      {stage045[92], stage045[93], stage045[94], stage045[95], stage045[96], stage045[97]},
      {stage047[60], stage047[61], stage047[62], stage047[63], stage047[64], stage047[65]},
      {stage049[138], stage048[146], stage047[148], stage046[160], stage045[198]}
   );
   gpc606_5 gpc606_5_1545(
      {stage045[98], stage045[99], stage045[100], stage045[101], stage045[102], stage045[103]},
      {stage047[66], stage047[67], stage047[68], stage047[69], stage047[70], stage047[71]},
      {stage049[139], stage048[147], stage047[149], stage046[161], stage045[199]}
   );
   gpc606_5 gpc606_5_1546(
      {stage045[104], stage045[105], stage045[106], stage045[107], stage045[108], stage045[109]},
      {stage047[72], stage047[73], stage047[74], stage047[75], stage047[76], stage047[77]},
      {stage049[140], stage048[148], stage047[150], stage046[162], stage045[200]}
   );
   gpc606_5 gpc606_5_1547(
      {stage045[110], stage045[111], stage045[112], stage045[113], stage045[114], stage045[115]},
      {stage047[78], stage047[79], stage047[80], stage047[81], stage047[82], stage047[83]},
      {stage049[141], stage048[149], stage047[151], stage046[163], stage045[201]}
   );
   gpc606_5 gpc606_5_1548(
      {stage045[116], stage045[117], stage045[118], stage045[119], stage045[120], stage045[121]},
      {stage047[84], stage047[85], stage047[86], stage047[87], stage047[88], stage047[89]},
      {stage049[142], stage048[150], stage047[152], stage046[164], stage045[202]}
   );
   gpc606_5 gpc606_5_1549(
      {stage045[122], stage045[123], stage045[124], stage045[125], stage045[126], stage045[127]},
      {stage047[90], stage047[91], stage047[92], stage047[93], stage047[94], stage047[95]},
      {stage049[143], stage048[151], stage047[153], stage046[165], stage045[203]}
   );
   gpc1_1 gpc1_1_1550(
      {stage046[50]},
      {stage046[166]}
   );
   gpc1_1 gpc1_1_1551(
      {stage046[51]},
      {stage046[167]}
   );
   gpc1_1 gpc1_1_1552(
      {stage046[52]},
      {stage046[168]}
   );
   gpc1_1 gpc1_1_1553(
      {stage046[53]},
      {stage046[169]}
   );
   gpc1_1 gpc1_1_1554(
      {stage046[54]},
      {stage046[170]}
   );
   gpc1_1 gpc1_1_1555(
      {stage046[55]},
      {stage046[171]}
   );
   gpc1_1 gpc1_1_1556(
      {stage046[56]},
      {stage046[172]}
   );
   gpc1_1 gpc1_1_1557(
      {stage046[57]},
      {stage046[173]}
   );
   gpc1_1 gpc1_1_1558(
      {stage046[58]},
      {stage046[174]}
   );
   gpc1_1 gpc1_1_1559(
      {stage046[59]},
      {stage046[175]}
   );
   gpc1_1 gpc1_1_1560(
      {stage046[60]},
      {stage046[176]}
   );
   gpc1_1 gpc1_1_1561(
      {stage046[61]},
      {stage046[177]}
   );
   gpc1_1 gpc1_1_1562(
      {stage046[62]},
      {stage046[178]}
   );
   gpc1_1 gpc1_1_1563(
      {stage046[63]},
      {stage046[179]}
   );
   gpc1_1 gpc1_1_1564(
      {stage046[64]},
      {stage046[180]}
   );
   gpc1_1 gpc1_1_1565(
      {stage046[65]},
      {stage046[181]}
   );
   gpc1_1 gpc1_1_1566(
      {stage046[66]},
      {stage046[182]}
   );
   gpc1_1 gpc1_1_1567(
      {stage046[67]},
      {stage046[183]}
   );
   gpc1_1 gpc1_1_1568(
      {stage046[68]},
      {stage046[184]}
   );
   gpc1_1 gpc1_1_1569(
      {stage046[69]},
      {stage046[185]}
   );
   gpc1_1 gpc1_1_1570(
      {stage046[70]},
      {stage046[186]}
   );
   gpc1_1 gpc1_1_1571(
      {stage046[71]},
      {stage046[187]}
   );
   gpc1_1 gpc1_1_1572(
      {stage046[72]},
      {stage046[188]}
   );
   gpc1_1 gpc1_1_1573(
      {stage046[73]},
      {stage046[189]}
   );
   gpc1_1 gpc1_1_1574(
      {stage046[74]},
      {stage046[190]}
   );
   gpc1_1 gpc1_1_1575(
      {stage046[75]},
      {stage046[191]}
   );
   gpc1_1 gpc1_1_1576(
      {stage046[76]},
      {stage046[192]}
   );
   gpc1_1 gpc1_1_1577(
      {stage046[77]},
      {stage046[193]}
   );
   gpc1_1 gpc1_1_1578(
      {stage046[78]},
      {stage046[194]}
   );
   gpc1_1 gpc1_1_1579(
      {stage046[79]},
      {stage046[195]}
   );
   gpc1_1 gpc1_1_1580(
      {stage046[80]},
      {stage046[196]}
   );
   gpc1_1 gpc1_1_1581(
      {stage046[81]},
      {stage046[197]}
   );
   gpc1_1 gpc1_1_1582(
      {stage046[82]},
      {stage046[198]}
   );
   gpc1_1 gpc1_1_1583(
      {stage046[83]},
      {stage046[199]}
   );
   gpc1_1 gpc1_1_1584(
      {stage046[84]},
      {stage046[200]}
   );
   gpc1_1 gpc1_1_1585(
      {stage046[85]},
      {stage046[201]}
   );
   gpc1_1 gpc1_1_1586(
      {stage046[86]},
      {stage046[202]}
   );
   gpc1_1 gpc1_1_1587(
      {stage046[87]},
      {stage046[203]}
   );
   gpc1_1 gpc1_1_1588(
      {stage046[88]},
      {stage046[204]}
   );
   gpc1_1 gpc1_1_1589(
      {stage046[89]},
      {stage046[205]}
   );
   gpc1_1 gpc1_1_1590(
      {stage046[90]},
      {stage046[206]}
   );
   gpc1_1 gpc1_1_1591(
      {stage046[91]},
      {stage046[207]}
   );
   gpc1_1 gpc1_1_1592(
      {stage046[92]},
      {stage046[208]}
   );
   gpc1_1 gpc1_1_1593(
      {stage046[93]},
      {stage046[209]}
   );
   gpc615_5 gpc615_5_1594(
      {stage046[94], stage046[95], stage046[96], stage046[97], stage046[98]},
      {stage047[96]},
      {stage048[0], stage048[1], stage048[2], stage048[3], stage048[4], stage048[5]},
      {stage050[128], stage049[144], stage048[152], stage047[154], stage046[210]}
   );
   gpc615_5 gpc615_5_1595(
      {stage046[99], stage046[100], stage046[101], stage046[102], stage046[103]},
      {stage047[97]},
      {stage048[6], stage048[7], stage048[8], stage048[9], stage048[10], stage048[11]},
      {stage050[129], stage049[145], stage048[153], stage047[155], stage046[211]}
   );
   gpc1406_5 gpc1406_5_1596(
      {stage046[104], stage046[105], stage046[106], stage046[107], stage046[108], stage046[109]},
      {stage048[12], stage048[13], stage048[14], stage048[15]},
      {stage049[0]},
      {stage050[130], stage049[146], stage048[154], stage047[156], stage046[212]}
   );
   gpc1406_5 gpc1406_5_1597(
      {stage046[110], stage046[111], stage046[112], stage046[113], stage046[114], stage046[115]},
      {stage048[16], stage048[17], stage048[18], stage048[19]},
      {stage049[1]},
      {stage050[131], stage049[147], stage048[155], stage047[157], stage046[213]}
   );
   gpc1406_5 gpc1406_5_1598(
      {stage046[116], stage046[117], stage046[118], stage046[119], stage046[120], stage046[121]},
      {stage048[20], stage048[21], stage048[22], stage048[23]},
      {stage049[2]},
      {stage050[132], stage049[148], stage048[156], stage047[158], stage046[214]}
   );
   gpc1406_5 gpc1406_5_1599(
      {stage046[122], stage046[123], stage046[124], stage046[125], stage046[126], stage046[127]},
      {stage048[24], stage048[25], stage048[26], stage048[27]},
      {stage049[3]},
      {stage050[133], stage049[149], stage048[157], stage047[159], stage046[215]}
   );
   gpc1_1 gpc1_1_1600(
      {stage047[98]},
      {stage047[160]}
   );
   gpc1_1 gpc1_1_1601(
      {stage047[99]},
      {stage047[161]}
   );
   gpc1_1 gpc1_1_1602(
      {stage047[100]},
      {stage047[162]}
   );
   gpc1_1 gpc1_1_1603(
      {stage047[101]},
      {stage047[163]}
   );
   gpc1_1 gpc1_1_1604(
      {stage047[102]},
      {stage047[164]}
   );
   gpc615_5 gpc615_5_1605(
      {stage047[103], stage047[104], stage047[105], stage047[106], stage047[107]},
      {stage048[28]},
      {stage049[4], stage049[5], stage049[6], stage049[7], stage049[8], stage049[9]},
      {stage051[128], stage050[134], stage049[150], stage048[158], stage047[165]}
   );
   gpc615_5 gpc615_5_1606(
      {stage047[108], stage047[109], stage047[110], stage047[111], stage047[112]},
      {stage048[29]},
      {stage049[10], stage049[11], stage049[12], stage049[13], stage049[14], stage049[15]},
      {stage051[129], stage050[135], stage049[151], stage048[159], stage047[166]}
   );
   gpc615_5 gpc615_5_1607(
      {stage047[113], stage047[114], stage047[115], stage047[116], stage047[117]},
      {stage048[30]},
      {stage049[16], stage049[17], stage049[18], stage049[19], stage049[20], stage049[21]},
      {stage051[130], stage050[136], stage049[152], stage048[160], stage047[167]}
   );
   gpc615_5 gpc615_5_1608(
      {stage047[118], stage047[119], stage047[120], stage047[121], stage047[122]},
      {stage048[31]},
      {stage049[22], stage049[23], stage049[24], stage049[25], stage049[26], stage049[27]},
      {stage051[131], stage050[137], stage049[153], stage048[161], stage047[168]}
   );
   gpc615_5 gpc615_5_1609(
      {stage047[123], stage047[124], stage047[125], stage047[126], stage047[127]},
      {stage048[32]},
      {stage049[28], stage049[29], stage049[30], stage049[31], stage049[32], stage049[33]},
      {stage051[132], stage050[138], stage049[154], stage048[162], stage047[169]}
   );
   gpc1_1 gpc1_1_1610(
      {stage048[33]},
      {stage048[163]}
   );
   gpc1_1 gpc1_1_1611(
      {stage048[34]},
      {stage048[164]}
   );
   gpc1_1 gpc1_1_1612(
      {stage048[35]},
      {stage048[165]}
   );
   gpc1_1 gpc1_1_1613(
      {stage048[36]},
      {stage048[166]}
   );
   gpc1_1 gpc1_1_1614(
      {stage048[37]},
      {stage048[167]}
   );
   gpc1_1 gpc1_1_1615(
      {stage048[38]},
      {stage048[168]}
   );
   gpc1_1 gpc1_1_1616(
      {stage048[39]},
      {stage048[169]}
   );
   gpc1_1 gpc1_1_1617(
      {stage048[40]},
      {stage048[170]}
   );
   gpc1_1 gpc1_1_1618(
      {stage048[41]},
      {stage048[171]}
   );
   gpc1_1 gpc1_1_1619(
      {stage048[42]},
      {stage048[172]}
   );
   gpc1_1 gpc1_1_1620(
      {stage048[43]},
      {stage048[173]}
   );
   gpc1_1 gpc1_1_1621(
      {stage048[44]},
      {stage048[174]}
   );
   gpc1_1 gpc1_1_1622(
      {stage048[45]},
      {stage048[175]}
   );
   gpc1_1 gpc1_1_1623(
      {stage048[46]},
      {stage048[176]}
   );
   gpc1_1 gpc1_1_1624(
      {stage048[47]},
      {stage048[177]}
   );
   gpc1_1 gpc1_1_1625(
      {stage048[48]},
      {stage048[178]}
   );
   gpc1_1 gpc1_1_1626(
      {stage048[49]},
      {stage048[179]}
   );
   gpc1_1 gpc1_1_1627(
      {stage048[50]},
      {stage048[180]}
   );
   gpc1_1 gpc1_1_1628(
      {stage048[51]},
      {stage048[181]}
   );
   gpc1_1 gpc1_1_1629(
      {stage048[52]},
      {stage048[182]}
   );
   gpc1_1 gpc1_1_1630(
      {stage048[53]},
      {stage048[183]}
   );
   gpc1_1 gpc1_1_1631(
      {stage048[54]},
      {stage048[184]}
   );
   gpc1_1 gpc1_1_1632(
      {stage048[55]},
      {stage048[185]}
   );
   gpc1_1 gpc1_1_1633(
      {stage048[56]},
      {stage048[186]}
   );
   gpc1_1 gpc1_1_1634(
      {stage048[57]},
      {stage048[187]}
   );
   gpc1_1 gpc1_1_1635(
      {stage048[58]},
      {stage048[188]}
   );
   gpc1_1 gpc1_1_1636(
      {stage048[59]},
      {stage048[189]}
   );
   gpc1_1 gpc1_1_1637(
      {stage048[60]},
      {stage048[190]}
   );
   gpc1_1 gpc1_1_1638(
      {stage048[61]},
      {stage048[191]}
   );
   gpc1_1 gpc1_1_1639(
      {stage048[62]},
      {stage048[192]}
   );
   gpc1_1 gpc1_1_1640(
      {stage048[63]},
      {stage048[193]}
   );
   gpc1_1 gpc1_1_1641(
      {stage048[64]},
      {stage048[194]}
   );
   gpc1_1 gpc1_1_1642(
      {stage048[65]},
      {stage048[195]}
   );
   gpc1_1 gpc1_1_1643(
      {stage048[66]},
      {stage048[196]}
   );
   gpc1_1 gpc1_1_1644(
      {stage048[67]},
      {stage048[197]}
   );
   gpc1_1 gpc1_1_1645(
      {stage048[68]},
      {stage048[198]}
   );
   gpc1_1 gpc1_1_1646(
      {stage048[69]},
      {stage048[199]}
   );
   gpc1_1 gpc1_1_1647(
      {stage048[70]},
      {stage048[200]}
   );
   gpc1_1 gpc1_1_1648(
      {stage048[71]},
      {stage048[201]}
   );
   gpc1_1 gpc1_1_1649(
      {stage048[72]},
      {stage048[202]}
   );
   gpc1_1 gpc1_1_1650(
      {stage048[73]},
      {stage048[203]}
   );
   gpc1_1 gpc1_1_1651(
      {stage048[74]},
      {stage048[204]}
   );
   gpc1_1 gpc1_1_1652(
      {stage048[75]},
      {stage048[205]}
   );
   gpc1_1 gpc1_1_1653(
      {stage048[76]},
      {stage048[206]}
   );
   gpc1_1 gpc1_1_1654(
      {stage048[77]},
      {stage048[207]}
   );
   gpc1_1 gpc1_1_1655(
      {stage048[78]},
      {stage048[208]}
   );
   gpc1_1 gpc1_1_1656(
      {stage048[79]},
      {stage048[209]}
   );
   gpc1_1 gpc1_1_1657(
      {stage048[80]},
      {stage048[210]}
   );
   gpc1_1 gpc1_1_1658(
      {stage048[81]},
      {stage048[211]}
   );
   gpc1_1 gpc1_1_1659(
      {stage048[82]},
      {stage048[212]}
   );
   gpc1_1 gpc1_1_1660(
      {stage048[83]},
      {stage048[213]}
   );
   gpc1_1 gpc1_1_1661(
      {stage048[84]},
      {stage048[214]}
   );
   gpc1_1 gpc1_1_1662(
      {stage048[85]},
      {stage048[215]}
   );
   gpc1_1 gpc1_1_1663(
      {stage048[86]},
      {stage048[216]}
   );
   gpc1_1 gpc1_1_1664(
      {stage048[87]},
      {stage048[217]}
   );
   gpc1_1 gpc1_1_1665(
      {stage048[88]},
      {stage048[218]}
   );
   gpc1_1 gpc1_1_1666(
      {stage048[89]},
      {stage048[219]}
   );
   gpc623_5 gpc623_5_1667(
      {stage048[90], stage048[91], stage048[92]},
      {stage049[34], stage049[35]},
      {stage050[0], stage050[1], stage050[2], stage050[3], stage050[4], stage050[5]},
      {stage052[128], stage051[133], stage050[139], stage049[155], stage048[220]}
   );
   gpc623_5 gpc623_5_1668(
      {stage048[93], stage048[94], stage048[95]},
      {stage049[36], stage049[37]},
      {stage050[6], stage050[7], stage050[8], stage050[9], stage050[10], stage050[11]},
      {stage052[129], stage051[134], stage050[140], stage049[156], stage048[221]}
   );
   gpc623_5 gpc623_5_1669(
      {stage048[96], stage048[97], stage048[98]},
      {stage049[38], stage049[39]},
      {stage050[12], stage050[13], stage050[14], stage050[15], stage050[16], stage050[17]},
      {stage052[130], stage051[135], stage050[141], stage049[157], stage048[222]}
   );
   gpc623_5 gpc623_5_1670(
      {stage048[99], stage048[100], stage048[101]},
      {stage049[40], stage049[41]},
      {stage050[18], stage050[19], stage050[20], stage050[21], stage050[22], stage050[23]},
      {stage052[131], stage051[136], stage050[142], stage049[158], stage048[223]}
   );
   gpc623_5 gpc623_5_1671(
      {stage048[102], stage048[103], stage048[104]},
      {stage049[42], stage049[43]},
      {stage050[24], stage050[25], stage050[26], stage050[27], stage050[28], stage050[29]},
      {stage052[132], stage051[137], stage050[143], stage049[159], stage048[224]}
   );
   gpc623_5 gpc623_5_1672(
      {stage048[105], stage048[106], stage048[107]},
      {stage049[44], stage049[45]},
      {stage050[30], stage050[31], stage050[32], stage050[33], stage050[34], stage050[35]},
      {stage052[133], stage051[138], stage050[144], stage049[160], stage048[225]}
   );
   gpc615_5 gpc615_5_1673(
      {stage048[108], stage048[109], stage048[110], stage048[111], stage048[112]},
      {stage049[46]},
      {stage050[36], stage050[37], stage050[38], stage050[39], stage050[40], stage050[41]},
      {stage052[134], stage051[139], stage050[145], stage049[161], stage048[226]}
   );
   gpc615_5 gpc615_5_1674(
      {stage048[113], stage048[114], stage048[115], stage048[116], stage048[117]},
      {stage049[47]},
      {stage050[42], stage050[43], stage050[44], stage050[45], stage050[46], stage050[47]},
      {stage052[135], stage051[140], stage050[146], stage049[162], stage048[227]}
   );
   gpc615_5 gpc615_5_1675(
      {stage048[118], stage048[119], stage048[120], stage048[121], stage048[122]},
      {stage049[48]},
      {stage050[48], stage050[49], stage050[50], stage050[51], stage050[52], stage050[53]},
      {stage052[136], stage051[141], stage050[147], stage049[163], stage048[228]}
   );
   gpc615_5 gpc615_5_1676(
      {stage048[123], stage048[124], stage048[125], stage048[126], stage048[127]},
      {stage049[49]},
      {stage050[54], stage050[55], stage050[56], stage050[57], stage050[58], stage050[59]},
      {stage052[137], stage051[142], stage050[148], stage049[164], stage048[229]}
   );
   gpc1_1 gpc1_1_1677(
      {stage049[50]},
      {stage049[165]}
   );
   gpc1_1 gpc1_1_1678(
      {stage049[51]},
      {stage049[166]}
   );
   gpc1_1 gpc1_1_1679(
      {stage049[52]},
      {stage049[167]}
   );
   gpc1_1 gpc1_1_1680(
      {stage049[53]},
      {stage049[168]}
   );
   gpc1_1 gpc1_1_1681(
      {stage049[54]},
      {stage049[169]}
   );
   gpc1_1 gpc1_1_1682(
      {stage049[55]},
      {stage049[170]}
   );
   gpc1_1 gpc1_1_1683(
      {stage049[56]},
      {stage049[171]}
   );
   gpc1_1 gpc1_1_1684(
      {stage049[57]},
      {stage049[172]}
   );
   gpc1_1 gpc1_1_1685(
      {stage049[58]},
      {stage049[173]}
   );
   gpc1_1 gpc1_1_1686(
      {stage049[59]},
      {stage049[174]}
   );
   gpc1_1 gpc1_1_1687(
      {stage049[60]},
      {stage049[175]}
   );
   gpc1_1 gpc1_1_1688(
      {stage049[61]},
      {stage049[176]}
   );
   gpc1_1 gpc1_1_1689(
      {stage049[62]},
      {stage049[177]}
   );
   gpc1_1 gpc1_1_1690(
      {stage049[63]},
      {stage049[178]}
   );
   gpc1_1 gpc1_1_1691(
      {stage049[64]},
      {stage049[179]}
   );
   gpc1_1 gpc1_1_1692(
      {stage049[65]},
      {stage049[180]}
   );
   gpc1_1 gpc1_1_1693(
      {stage049[66]},
      {stage049[181]}
   );
   gpc1_1 gpc1_1_1694(
      {stage049[67]},
      {stage049[182]}
   );
   gpc1_1 gpc1_1_1695(
      {stage049[68]},
      {stage049[183]}
   );
   gpc1_1 gpc1_1_1696(
      {stage049[69]},
      {stage049[184]}
   );
   gpc1_1 gpc1_1_1697(
      {stage049[70]},
      {stage049[185]}
   );
   gpc1_1 gpc1_1_1698(
      {stage049[71]},
      {stage049[186]}
   );
   gpc1_1 gpc1_1_1699(
      {stage049[72]},
      {stage049[187]}
   );
   gpc1_1 gpc1_1_1700(
      {stage049[73]},
      {stage049[188]}
   );
   gpc1_1 gpc1_1_1701(
      {stage049[74]},
      {stage049[189]}
   );
   gpc1_1 gpc1_1_1702(
      {stage049[75]},
      {stage049[190]}
   );
   gpc1_1 gpc1_1_1703(
      {stage049[76]},
      {stage049[191]}
   );
   gpc1_1 gpc1_1_1704(
      {stage049[77]},
      {stage049[192]}
   );
   gpc1_1 gpc1_1_1705(
      {stage049[78]},
      {stage049[193]}
   );
   gpc1_1 gpc1_1_1706(
      {stage049[79]},
      {stage049[194]}
   );
   gpc1_1 gpc1_1_1707(
      {stage049[80]},
      {stage049[195]}
   );
   gpc606_5 gpc606_5_1708(
      {stage049[81], stage049[82], stage049[83], stage049[84], stage049[85], stage049[86]},
      {stage051[0], stage051[1], stage051[2], stage051[3], stage051[4], stage051[5]},
      {stage053[128], stage052[138], stage051[143], stage050[149], stage049[196]}
   );
   gpc606_5 gpc606_5_1709(
      {stage049[87], stage049[88], stage049[89], stage049[90], stage049[91], stage049[92]},
      {stage051[6], stage051[7], stage051[8], stage051[9], stage051[10], stage051[11]},
      {stage053[129], stage052[139], stage051[144], stage050[150], stage049[197]}
   );
   gpc606_5 gpc606_5_1710(
      {stage049[93], stage049[94], stage049[95], stage049[96], stage049[97], stage049[98]},
      {stage051[12], stage051[13], stage051[14], stage051[15], stage051[16], stage051[17]},
      {stage053[130], stage052[140], stage051[145], stage050[151], stage049[198]}
   );
   gpc606_5 gpc606_5_1711(
      {stage049[99], stage049[100], stage049[101], stage049[102], stage049[103], stage049[104]},
      {stage051[18], stage051[19], stage051[20], stage051[21], stage051[22], stage051[23]},
      {stage053[131], stage052[141], stage051[146], stage050[152], stage049[199]}
   );
   gpc606_5 gpc606_5_1712(
      {stage049[105], stage049[106], stage049[107], stage049[108], stage049[109], stage049[110]},
      {stage051[24], stage051[25], stage051[26], stage051[27], stage051[28], stage051[29]},
      {stage053[132], stage052[142], stage051[147], stage050[153], stage049[200]}
   );
   gpc606_5 gpc606_5_1713(
      {stage049[111], stage049[112], stage049[113], stage049[114], stage049[115], stage049[116]},
      {stage051[30], stage051[31], stage051[32], stage051[33], stage051[34], stage051[35]},
      {stage053[133], stage052[143], stage051[148], stage050[154], stage049[201]}
   );
   gpc606_5 gpc606_5_1714(
      {stage049[117], stage049[118], stage049[119], stage049[120], stage049[121], stage049[122]},
      {stage051[36], stage051[37], stage051[38], stage051[39], stage051[40], stage051[41]},
      {stage053[134], stage052[144], stage051[149], stage050[155], stage049[202]}
   );
   gpc615_5 gpc615_5_1715(
      {stage049[123], stage049[124], stage049[125], stage049[126], stage049[127]},
      {stage050[60]},
      {stage051[42], stage051[43], stage051[44], stage051[45], stage051[46], stage051[47]},
      {stage053[135], stage052[145], stage051[150], stage050[156], stage049[203]}
   );
   gpc1_1 gpc1_1_1716(
      {stage050[61]},
      {stage050[157]}
   );
   gpc1_1 gpc1_1_1717(
      {stage050[62]},
      {stage050[158]}
   );
   gpc1_1 gpc1_1_1718(
      {stage050[63]},
      {stage050[159]}
   );
   gpc1_1 gpc1_1_1719(
      {stage050[64]},
      {stage050[160]}
   );
   gpc1_1 gpc1_1_1720(
      {stage050[65]},
      {stage050[161]}
   );
   gpc1_1 gpc1_1_1721(
      {stage050[66]},
      {stage050[162]}
   );
   gpc1_1 gpc1_1_1722(
      {stage050[67]},
      {stage050[163]}
   );
   gpc1_1 gpc1_1_1723(
      {stage050[68]},
      {stage050[164]}
   );
   gpc1_1 gpc1_1_1724(
      {stage050[69]},
      {stage050[165]}
   );
   gpc1_1 gpc1_1_1725(
      {stage050[70]},
      {stage050[166]}
   );
   gpc1_1 gpc1_1_1726(
      {stage050[71]},
      {stage050[167]}
   );
   gpc1_1 gpc1_1_1727(
      {stage050[72]},
      {stage050[168]}
   );
   gpc1_1 gpc1_1_1728(
      {stage050[73]},
      {stage050[169]}
   );
   gpc1_1 gpc1_1_1729(
      {stage050[74]},
      {stage050[170]}
   );
   gpc1_1 gpc1_1_1730(
      {stage050[75]},
      {stage050[171]}
   );
   gpc1_1 gpc1_1_1731(
      {stage050[76]},
      {stage050[172]}
   );
   gpc1_1 gpc1_1_1732(
      {stage050[77]},
      {stage050[173]}
   );
   gpc1_1 gpc1_1_1733(
      {stage050[78]},
      {stage050[174]}
   );
   gpc1_1 gpc1_1_1734(
      {stage050[79]},
      {stage050[175]}
   );
   gpc1_1 gpc1_1_1735(
      {stage050[80]},
      {stage050[176]}
   );
   gpc1_1 gpc1_1_1736(
      {stage050[81]},
      {stage050[177]}
   );
   gpc1_1 gpc1_1_1737(
      {stage050[82]},
      {stage050[178]}
   );
   gpc1_1 gpc1_1_1738(
      {stage050[83]},
      {stage050[179]}
   );
   gpc1_1 gpc1_1_1739(
      {stage050[84]},
      {stage050[180]}
   );
   gpc1_1 gpc1_1_1740(
      {stage050[85]},
      {stage050[181]}
   );
   gpc1_1 gpc1_1_1741(
      {stage050[86]},
      {stage050[182]}
   );
   gpc1_1 gpc1_1_1742(
      {stage050[87]},
      {stage050[183]}
   );
   gpc1_1 gpc1_1_1743(
      {stage050[88]},
      {stage050[184]}
   );
   gpc1_1 gpc1_1_1744(
      {stage050[89]},
      {stage050[185]}
   );
   gpc1_1 gpc1_1_1745(
      {stage050[90]},
      {stage050[186]}
   );
   gpc1_1 gpc1_1_1746(
      {stage050[91]},
      {stage050[187]}
   );
   gpc1_1 gpc1_1_1747(
      {stage050[92]},
      {stage050[188]}
   );
   gpc1_1 gpc1_1_1748(
      {stage050[93]},
      {stage050[189]}
   );
   gpc1_1 gpc1_1_1749(
      {stage050[94]},
      {stage050[190]}
   );
   gpc1_1 gpc1_1_1750(
      {stage050[95]},
      {stage050[191]}
   );
   gpc1_1 gpc1_1_1751(
      {stage050[96]},
      {stage050[192]}
   );
   gpc1_1 gpc1_1_1752(
      {stage050[97]},
      {stage050[193]}
   );
   gpc1_1 gpc1_1_1753(
      {stage050[98]},
      {stage050[194]}
   );
   gpc1_1 gpc1_1_1754(
      {stage050[99]},
      {stage050[195]}
   );
   gpc1_1 gpc1_1_1755(
      {stage050[100]},
      {stage050[196]}
   );
   gpc1_1 gpc1_1_1756(
      {stage050[101]},
      {stage050[197]}
   );
   gpc1_1 gpc1_1_1757(
      {stage050[102]},
      {stage050[198]}
   );
   gpc1_1 gpc1_1_1758(
      {stage050[103]},
      {stage050[199]}
   );
   gpc1_1 gpc1_1_1759(
      {stage050[104]},
      {stage050[200]}
   );
   gpc1_1 gpc1_1_1760(
      {stage050[105]},
      {stage050[201]}
   );
   gpc1_1 gpc1_1_1761(
      {stage050[106]},
      {stage050[202]}
   );
   gpc1_1 gpc1_1_1762(
      {stage050[107]},
      {stage050[203]}
   );
   gpc1_1 gpc1_1_1763(
      {stage050[108]},
      {stage050[204]}
   );
   gpc1_1 gpc1_1_1764(
      {stage050[109]},
      {stage050[205]}
   );
   gpc1_1 gpc1_1_1765(
      {stage050[110]},
      {stage050[206]}
   );
   gpc1_1 gpc1_1_1766(
      {stage050[111]},
      {stage050[207]}
   );
   gpc1_1 gpc1_1_1767(
      {stage050[112]},
      {stage050[208]}
   );
   gpc1_1 gpc1_1_1768(
      {stage050[113]},
      {stage050[209]}
   );
   gpc1_1 gpc1_1_1769(
      {stage050[114]},
      {stage050[210]}
   );
   gpc1_1 gpc1_1_1770(
      {stage050[115]},
      {stage050[211]}
   );
   gpc1_1 gpc1_1_1771(
      {stage050[116]},
      {stage050[212]}
   );
   gpc1_1 gpc1_1_1772(
      {stage050[117]},
      {stage050[213]}
   );
   gpc1_1 gpc1_1_1773(
      {stage050[118]},
      {stage050[214]}
   );
   gpc1_1 gpc1_1_1774(
      {stage050[119]},
      {stage050[215]}
   );
   gpc1_1 gpc1_1_1775(
      {stage050[120]},
      {stage050[216]}
   );
   gpc1_1 gpc1_1_1776(
      {stage050[121]},
      {stage050[217]}
   );
   gpc1_1 gpc1_1_1777(
      {stage050[122]},
      {stage050[218]}
   );
   gpc1_1 gpc1_1_1778(
      {stage050[123]},
      {stage050[219]}
   );
   gpc1_1 gpc1_1_1779(
      {stage050[124]},
      {stage050[220]}
   );
   gpc1_1 gpc1_1_1780(
      {stage050[125]},
      {stage050[221]}
   );
   gpc1_1 gpc1_1_1781(
      {stage050[126]},
      {stage050[222]}
   );
   gpc1_1 gpc1_1_1782(
      {stage050[127]},
      {stage050[223]}
   );
   gpc615_5 gpc615_5_1783(
      {stage051[48], stage051[49], stage051[50], stage051[51], stage051[52]},
      {stage052[0]},
      {stage053[0], stage053[1], stage053[2], stage053[3], stage053[4], stage053[5]},
      {stage055[128], stage054[128], stage053[136], stage052[146], stage051[151]}
   );
   gpc615_5 gpc615_5_1784(
      {stage051[53], stage051[54], stage051[55], stage051[56], stage051[57]},
      {stage052[1]},
      {stage053[6], stage053[7], stage053[8], stage053[9], stage053[10], stage053[11]},
      {stage055[129], stage054[129], stage053[137], stage052[147], stage051[152]}
   );
   gpc615_5 gpc615_5_1785(
      {stage051[58], stage051[59], stage051[60], stage051[61], stage051[62]},
      {stage052[2]},
      {stage053[12], stage053[13], stage053[14], stage053[15], stage053[16], stage053[17]},
      {stage055[130], stage054[130], stage053[138], stage052[148], stage051[153]}
   );
   gpc615_5 gpc615_5_1786(
      {stage051[63], stage051[64], stage051[65], stage051[66], stage051[67]},
      {stage052[3]},
      {stage053[18], stage053[19], stage053[20], stage053[21], stage053[22], stage053[23]},
      {stage055[131], stage054[131], stage053[139], stage052[149], stage051[154]}
   );
   gpc615_5 gpc615_5_1787(
      {stage051[68], stage051[69], stage051[70], stage051[71], stage051[72]},
      {stage052[4]},
      {stage053[24], stage053[25], stage053[26], stage053[27], stage053[28], stage053[29]},
      {stage055[132], stage054[132], stage053[140], stage052[150], stage051[155]}
   );
   gpc615_5 gpc615_5_1788(
      {stage051[73], stage051[74], stage051[75], stage051[76], stage051[77]},
      {stage052[5]},
      {stage053[30], stage053[31], stage053[32], stage053[33], stage053[34], stage053[35]},
      {stage055[133], stage054[133], stage053[141], stage052[151], stage051[156]}
   );
   gpc615_5 gpc615_5_1789(
      {stage051[78], stage051[79], stage051[80], stage051[81], stage051[82]},
      {stage052[6]},
      {stage053[36], stage053[37], stage053[38], stage053[39], stage053[40], stage053[41]},
      {stage055[134], stage054[134], stage053[142], stage052[152], stage051[157]}
   );
   gpc615_5 gpc615_5_1790(
      {stage051[83], stage051[84], stage051[85], stage051[86], stage051[87]},
      {stage052[7]},
      {stage053[42], stage053[43], stage053[44], stage053[45], stage053[46], stage053[47]},
      {stage055[135], stage054[135], stage053[143], stage052[153], stage051[158]}
   );
   gpc615_5 gpc615_5_1791(
      {stage051[88], stage051[89], stage051[90], stage051[91], stage051[92]},
      {stage052[8]},
      {stage053[48], stage053[49], stage053[50], stage053[51], stage053[52], stage053[53]},
      {stage055[136], stage054[136], stage053[144], stage052[154], stage051[159]}
   );
   gpc615_5 gpc615_5_1792(
      {stage051[93], stage051[94], stage051[95], stage051[96], stage051[97]},
      {stage052[9]},
      {stage053[54], stage053[55], stage053[56], stage053[57], stage053[58], stage053[59]},
      {stage055[137], stage054[137], stage053[145], stage052[155], stage051[160]}
   );
   gpc615_5 gpc615_5_1793(
      {stage051[98], stage051[99], stage051[100], stage051[101], stage051[102]},
      {stage052[10]},
      {stage053[60], stage053[61], stage053[62], stage053[63], stage053[64], stage053[65]},
      {stage055[138], stage054[138], stage053[146], stage052[156], stage051[161]}
   );
   gpc615_5 gpc615_5_1794(
      {stage051[103], stage051[104], stage051[105], stage051[106], stage051[107]},
      {stage052[11]},
      {stage053[66], stage053[67], stage053[68], stage053[69], stage053[70], stage053[71]},
      {stage055[139], stage054[139], stage053[147], stage052[157], stage051[162]}
   );
   gpc615_5 gpc615_5_1795(
      {stage051[108], stage051[109], stage051[110], stage051[111], stage051[112]},
      {stage052[12]},
      {stage053[72], stage053[73], stage053[74], stage053[75], stage053[76], stage053[77]},
      {stage055[140], stage054[140], stage053[148], stage052[158], stage051[163]}
   );
   gpc615_5 gpc615_5_1796(
      {stage051[113], stage051[114], stage051[115], stage051[116], stage051[117]},
      {stage052[13]},
      {stage053[78], stage053[79], stage053[80], stage053[81], stage053[82], stage053[83]},
      {stage055[141], stage054[141], stage053[149], stage052[159], stage051[164]}
   );
   gpc615_5 gpc615_5_1797(
      {stage051[118], stage051[119], stage051[120], stage051[121], stage051[122]},
      {stage052[14]},
      {stage053[84], stage053[85], stage053[86], stage053[87], stage053[88], stage053[89]},
      {stage055[142], stage054[142], stage053[150], stage052[160], stage051[165]}
   );
   gpc615_5 gpc615_5_1798(
      {stage051[123], stage051[124], stage051[125], stage051[126], stage051[127]},
      {stage052[15]},
      {stage053[90], stage053[91], stage053[92], stage053[93], stage053[94], stage053[95]},
      {stage055[143], stage054[143], stage053[151], stage052[161], stage051[166]}
   );
   gpc1_1 gpc1_1_1799(
      {stage052[16]},
      {stage052[162]}
   );
   gpc1_1 gpc1_1_1800(
      {stage052[17]},
      {stage052[163]}
   );
   gpc1_1 gpc1_1_1801(
      {stage052[18]},
      {stage052[164]}
   );
   gpc1_1 gpc1_1_1802(
      {stage052[19]},
      {stage052[165]}
   );
   gpc1_1 gpc1_1_1803(
      {stage052[20]},
      {stage052[166]}
   );
   gpc1_1 gpc1_1_1804(
      {stage052[21]},
      {stage052[167]}
   );
   gpc1_1 gpc1_1_1805(
      {stage052[22]},
      {stage052[168]}
   );
   gpc1_1 gpc1_1_1806(
      {stage052[23]},
      {stage052[169]}
   );
   gpc1_1 gpc1_1_1807(
      {stage052[24]},
      {stage052[170]}
   );
   gpc1_1 gpc1_1_1808(
      {stage052[25]},
      {stage052[171]}
   );
   gpc1_1 gpc1_1_1809(
      {stage052[26]},
      {stage052[172]}
   );
   gpc1_1 gpc1_1_1810(
      {stage052[27]},
      {stage052[173]}
   );
   gpc1_1 gpc1_1_1811(
      {stage052[28]},
      {stage052[174]}
   );
   gpc1_1 gpc1_1_1812(
      {stage052[29]},
      {stage052[175]}
   );
   gpc1_1 gpc1_1_1813(
      {stage052[30]},
      {stage052[176]}
   );
   gpc1_1 gpc1_1_1814(
      {stage052[31]},
      {stage052[177]}
   );
   gpc1_1 gpc1_1_1815(
      {stage052[32]},
      {stage052[178]}
   );
   gpc1_1 gpc1_1_1816(
      {stage052[33]},
      {stage052[179]}
   );
   gpc1_1 gpc1_1_1817(
      {stage052[34]},
      {stage052[180]}
   );
   gpc1_1 gpc1_1_1818(
      {stage052[35]},
      {stage052[181]}
   );
   gpc1_1 gpc1_1_1819(
      {stage052[36]},
      {stage052[182]}
   );
   gpc1_1 gpc1_1_1820(
      {stage052[37]},
      {stage052[183]}
   );
   gpc1_1 gpc1_1_1821(
      {stage052[38]},
      {stage052[184]}
   );
   gpc1_1 gpc1_1_1822(
      {stage052[39]},
      {stage052[185]}
   );
   gpc1_1 gpc1_1_1823(
      {stage052[40]},
      {stage052[186]}
   );
   gpc1_1 gpc1_1_1824(
      {stage052[41]},
      {stage052[187]}
   );
   gpc1_1 gpc1_1_1825(
      {stage052[42]},
      {stage052[188]}
   );
   gpc1_1 gpc1_1_1826(
      {stage052[43]},
      {stage052[189]}
   );
   gpc1_1 gpc1_1_1827(
      {stage052[44]},
      {stage052[190]}
   );
   gpc1_1 gpc1_1_1828(
      {stage052[45]},
      {stage052[191]}
   );
   gpc1_1 gpc1_1_1829(
      {stage052[46]},
      {stage052[192]}
   );
   gpc1_1 gpc1_1_1830(
      {stage052[47]},
      {stage052[193]}
   );
   gpc1_1 gpc1_1_1831(
      {stage052[48]},
      {stage052[194]}
   );
   gpc1_1 gpc1_1_1832(
      {stage052[49]},
      {stage052[195]}
   );
   gpc1_1 gpc1_1_1833(
      {stage052[50]},
      {stage052[196]}
   );
   gpc1_1 gpc1_1_1834(
      {stage052[51]},
      {stage052[197]}
   );
   gpc1_1 gpc1_1_1835(
      {stage052[52]},
      {stage052[198]}
   );
   gpc1_1 gpc1_1_1836(
      {stage052[53]},
      {stage052[199]}
   );
   gpc1_1 gpc1_1_1837(
      {stage052[54]},
      {stage052[200]}
   );
   gpc1_1 gpc1_1_1838(
      {stage052[55]},
      {stage052[201]}
   );
   gpc606_5 gpc606_5_1839(
      {stage052[56], stage052[57], stage052[58], stage052[59], stage052[60], stage052[61]},
      {stage054[0], stage054[1], stage054[2], stage054[3], stage054[4], stage054[5]},
      {stage056[128], stage055[144], stage054[144], stage053[152], stage052[202]}
   );
   gpc606_5 gpc606_5_1840(
      {stage052[62], stage052[63], stage052[64], stage052[65], stage052[66], stage052[67]},
      {stage054[6], stage054[7], stage054[8], stage054[9], stage054[10], stage054[11]},
      {stage056[129], stage055[145], stage054[145], stage053[153], stage052[203]}
   );
   gpc606_5 gpc606_5_1841(
      {stage052[68], stage052[69], stage052[70], stage052[71], stage052[72], stage052[73]},
      {stage054[12], stage054[13], stage054[14], stage054[15], stage054[16], stage054[17]},
      {stage056[130], stage055[146], stage054[146], stage053[154], stage052[204]}
   );
   gpc606_5 gpc606_5_1842(
      {stage052[74], stage052[75], stage052[76], stage052[77], stage052[78], stage052[79]},
      {stage054[18], stage054[19], stage054[20], stage054[21], stage054[22], stage054[23]},
      {stage056[131], stage055[147], stage054[147], stage053[155], stage052[205]}
   );
   gpc606_5 gpc606_5_1843(
      {stage052[80], stage052[81], stage052[82], stage052[83], stage052[84], stage052[85]},
      {stage054[24], stage054[25], stage054[26], stage054[27], stage054[28], stage054[29]},
      {stage056[132], stage055[148], stage054[148], stage053[156], stage052[206]}
   );
   gpc606_5 gpc606_5_1844(
      {stage052[86], stage052[87], stage052[88], stage052[89], stage052[90], stage052[91]},
      {stage054[30], stage054[31], stage054[32], stage054[33], stage054[34], stage054[35]},
      {stage056[133], stage055[149], stage054[149], stage053[157], stage052[207]}
   );
   gpc606_5 gpc606_5_1845(
      {stage052[92], stage052[93], stage052[94], stage052[95], stage052[96], stage052[97]},
      {stage054[36], stage054[37], stage054[38], stage054[39], stage054[40], stage054[41]},
      {stage056[134], stage055[150], stage054[150], stage053[158], stage052[208]}
   );
   gpc606_5 gpc606_5_1846(
      {stage052[98], stage052[99], stage052[100], stage052[101], stage052[102], stage052[103]},
      {stage054[42], stage054[43], stage054[44], stage054[45], stage054[46], stage054[47]},
      {stage056[135], stage055[151], stage054[151], stage053[159], stage052[209]}
   );
   gpc606_5 gpc606_5_1847(
      {stage052[104], stage052[105], stage052[106], stage052[107], stage052[108], stage052[109]},
      {stage054[48], stage054[49], stage054[50], stage054[51], stage054[52], stage054[53]},
      {stage056[136], stage055[152], stage054[152], stage053[160], stage052[210]}
   );
   gpc606_5 gpc606_5_1848(
      {stage052[110], stage052[111], stage052[112], stage052[113], stage052[114], stage052[115]},
      {stage054[54], stage054[55], stage054[56], stage054[57], stage054[58], stage054[59]},
      {stage056[137], stage055[153], stage054[153], stage053[161], stage052[211]}
   );
   gpc606_5 gpc606_5_1849(
      {stage052[116], stage052[117], stage052[118], stage052[119], stage052[120], stage052[121]},
      {stage054[60], stage054[61], stage054[62], stage054[63], stage054[64], stage054[65]},
      {stage056[138], stage055[154], stage054[154], stage053[162], stage052[212]}
   );
   gpc606_5 gpc606_5_1850(
      {stage052[122], stage052[123], stage052[124], stage052[125], stage052[126], stage052[127]},
      {stage054[66], stage054[67], stage054[68], stage054[69], stage054[70], stage054[71]},
      {stage056[139], stage055[155], stage054[155], stage053[163], stage052[213]}
   );
   gpc1_1 gpc1_1_1851(
      {stage053[96]},
      {stage053[164]}
   );
   gpc1_1 gpc1_1_1852(
      {stage053[97]},
      {stage053[165]}
   );
   gpc606_5 gpc606_5_1853(
      {stage053[98], stage053[99], stage053[100], stage053[101], stage053[102], stage053[103]},
      {stage055[0], stage055[1], stage055[2], stage055[3], stage055[4], stage055[5]},
      {stage057[128], stage056[140], stage055[156], stage054[156], stage053[166]}
   );
   gpc606_5 gpc606_5_1854(
      {stage053[104], stage053[105], stage053[106], stage053[107], stage053[108], stage053[109]},
      {stage055[6], stage055[7], stage055[8], stage055[9], stage055[10], stage055[11]},
      {stage057[129], stage056[141], stage055[157], stage054[157], stage053[167]}
   );
   gpc606_5 gpc606_5_1855(
      {stage053[110], stage053[111], stage053[112], stage053[113], stage053[114], stage053[115]},
      {stage055[12], stage055[13], stage055[14], stage055[15], stage055[16], stage055[17]},
      {stage057[130], stage056[142], stage055[158], stage054[158], stage053[168]}
   );
   gpc606_5 gpc606_5_1856(
      {stage053[116], stage053[117], stage053[118], stage053[119], stage053[120], stage053[121]},
      {stage055[18], stage055[19], stage055[20], stage055[21], stage055[22], stage055[23]},
      {stage057[131], stage056[143], stage055[159], stage054[159], stage053[169]}
   );
   gpc606_5 gpc606_5_1857(
      {stage053[122], stage053[123], stage053[124], stage053[125], stage053[126], stage053[127]},
      {stage055[24], stage055[25], stage055[26], stage055[27], stage055[28], stage055[29]},
      {stage057[132], stage056[144], stage055[160], stage054[160], stage053[170]}
   );
   gpc1_1 gpc1_1_1858(
      {stage054[72]},
      {stage054[161]}
   );
   gpc1_1 gpc1_1_1859(
      {stage054[73]},
      {stage054[162]}
   );
   gpc1_1 gpc1_1_1860(
      {stage054[74]},
      {stage054[163]}
   );
   gpc1_1 gpc1_1_1861(
      {stage054[75]},
      {stage054[164]}
   );
   gpc1_1 gpc1_1_1862(
      {stage054[76]},
      {stage054[165]}
   );
   gpc1_1 gpc1_1_1863(
      {stage054[77]},
      {stage054[166]}
   );
   gpc1_1 gpc1_1_1864(
      {stage054[78]},
      {stage054[167]}
   );
   gpc1_1 gpc1_1_1865(
      {stage054[79]},
      {stage054[168]}
   );
   gpc1_1 gpc1_1_1866(
      {stage054[80]},
      {stage054[169]}
   );
   gpc1_1 gpc1_1_1867(
      {stage054[81]},
      {stage054[170]}
   );
   gpc1_1 gpc1_1_1868(
      {stage054[82]},
      {stage054[171]}
   );
   gpc1_1 gpc1_1_1869(
      {stage054[83]},
      {stage054[172]}
   );
   gpc1_1 gpc1_1_1870(
      {stage054[84]},
      {stage054[173]}
   );
   gpc1_1 gpc1_1_1871(
      {stage054[85]},
      {stage054[174]}
   );
   gpc1_1 gpc1_1_1872(
      {stage054[86]},
      {stage054[175]}
   );
   gpc1_1 gpc1_1_1873(
      {stage054[87]},
      {stage054[176]}
   );
   gpc1_1 gpc1_1_1874(
      {stage054[88]},
      {stage054[177]}
   );
   gpc1_1 gpc1_1_1875(
      {stage054[89]},
      {stage054[178]}
   );
   gpc1_1 gpc1_1_1876(
      {stage054[90]},
      {stage054[179]}
   );
   gpc1_1 gpc1_1_1877(
      {stage054[91]},
      {stage054[180]}
   );
   gpc1_1 gpc1_1_1878(
      {stage054[92]},
      {stage054[181]}
   );
   gpc1_1 gpc1_1_1879(
      {stage054[93]},
      {stage054[182]}
   );
   gpc1_1 gpc1_1_1880(
      {stage054[94]},
      {stage054[183]}
   );
   gpc1_1 gpc1_1_1881(
      {stage054[95]},
      {stage054[184]}
   );
   gpc1_1 gpc1_1_1882(
      {stage054[96]},
      {stage054[185]}
   );
   gpc1_1 gpc1_1_1883(
      {stage054[97]},
      {stage054[186]}
   );
   gpc1_1 gpc1_1_1884(
      {stage054[98]},
      {stage054[187]}
   );
   gpc1_1 gpc1_1_1885(
      {stage054[99]},
      {stage054[188]}
   );
   gpc1_1 gpc1_1_1886(
      {stage054[100]},
      {stage054[189]}
   );
   gpc1_1 gpc1_1_1887(
      {stage054[101]},
      {stage054[190]}
   );
   gpc1_1 gpc1_1_1888(
      {stage054[102]},
      {stage054[191]}
   );
   gpc1_1 gpc1_1_1889(
      {stage054[103]},
      {stage054[192]}
   );
   gpc1_1 gpc1_1_1890(
      {stage054[104]},
      {stage054[193]}
   );
   gpc1_1 gpc1_1_1891(
      {stage054[105]},
      {stage054[194]}
   );
   gpc1_1 gpc1_1_1892(
      {stage054[106]},
      {stage054[195]}
   );
   gpc1_1 gpc1_1_1893(
      {stage054[107]},
      {stage054[196]}
   );
   gpc1_1 gpc1_1_1894(
      {stage054[108]},
      {stage054[197]}
   );
   gpc1_1 gpc1_1_1895(
      {stage054[109]},
      {stage054[198]}
   );
   gpc1_1 gpc1_1_1896(
      {stage054[110]},
      {stage054[199]}
   );
   gpc1_1 gpc1_1_1897(
      {stage054[111]},
      {stage054[200]}
   );
   gpc1_1 gpc1_1_1898(
      {stage054[112]},
      {stage054[201]}
   );
   gpc615_5 gpc615_5_1899(
      {stage054[113], stage054[114], stage054[115], stage054[116], stage054[117]},
      {stage055[30]},
      {stage056[0], stage056[1], stage056[2], stage056[3], stage056[4], stage056[5]},
      {stage058[128], stage057[133], stage056[145], stage055[161], stage054[202]}
   );
   gpc615_5 gpc615_5_1900(
      {stage054[118], stage054[119], stage054[120], stage054[121], stage054[122]},
      {stage055[31]},
      {stage056[6], stage056[7], stage056[8], stage056[9], stage056[10], stage056[11]},
      {stage058[129], stage057[134], stage056[146], stage055[162], stage054[203]}
   );
   gpc615_5 gpc615_5_1901(
      {stage054[123], stage054[124], stage054[125], stage054[126], stage054[127]},
      {stage055[32]},
      {stage056[12], stage056[13], stage056[14], stage056[15], stage056[16], stage056[17]},
      {stage058[130], stage057[135], stage056[147], stage055[163], stage054[204]}
   );
   gpc1_1 gpc1_1_1902(
      {stage055[33]},
      {stage055[164]}
   );
   gpc1_1 gpc1_1_1903(
      {stage055[34]},
      {stage055[165]}
   );
   gpc1_1 gpc1_1_1904(
      {stage055[35]},
      {stage055[166]}
   );
   gpc1_1 gpc1_1_1905(
      {stage055[36]},
      {stage055[167]}
   );
   gpc1_1 gpc1_1_1906(
      {stage055[37]},
      {stage055[168]}
   );
   gpc1_1 gpc1_1_1907(
      {stage055[38]},
      {stage055[169]}
   );
   gpc1_1 gpc1_1_1908(
      {stage055[39]},
      {stage055[170]}
   );
   gpc1_1 gpc1_1_1909(
      {stage055[40]},
      {stage055[171]}
   );
   gpc1_1 gpc1_1_1910(
      {stage055[41]},
      {stage055[172]}
   );
   gpc1_1 gpc1_1_1911(
      {stage055[42]},
      {stage055[173]}
   );
   gpc1_1 gpc1_1_1912(
      {stage055[43]},
      {stage055[174]}
   );
   gpc1_1 gpc1_1_1913(
      {stage055[44]},
      {stage055[175]}
   );
   gpc1_1 gpc1_1_1914(
      {stage055[45]},
      {stage055[176]}
   );
   gpc1_1 gpc1_1_1915(
      {stage055[46]},
      {stage055[177]}
   );
   gpc1_1 gpc1_1_1916(
      {stage055[47]},
      {stage055[178]}
   );
   gpc1_1 gpc1_1_1917(
      {stage055[48]},
      {stage055[179]}
   );
   gpc1_1 gpc1_1_1918(
      {stage055[49]},
      {stage055[180]}
   );
   gpc1_1 gpc1_1_1919(
      {stage055[50]},
      {stage055[181]}
   );
   gpc1_1 gpc1_1_1920(
      {stage055[51]},
      {stage055[182]}
   );
   gpc1_1 gpc1_1_1921(
      {stage055[52]},
      {stage055[183]}
   );
   gpc1_1 gpc1_1_1922(
      {stage055[53]},
      {stage055[184]}
   );
   gpc1_1 gpc1_1_1923(
      {stage055[54]},
      {stage055[185]}
   );
   gpc1_1 gpc1_1_1924(
      {stage055[55]},
      {stage055[186]}
   );
   gpc606_5 gpc606_5_1925(
      {stage055[56], stage055[57], stage055[58], stage055[59], stage055[60], stage055[61]},
      {stage057[0], stage057[1], stage057[2], stage057[3], stage057[4], stage057[5]},
      {stage059[128], stage058[131], stage057[136], stage056[148], stage055[187]}
   );
   gpc606_5 gpc606_5_1926(
      {stage055[62], stage055[63], stage055[64], stage055[65], stage055[66], stage055[67]},
      {stage057[6], stage057[7], stage057[8], stage057[9], stage057[10], stage057[11]},
      {stage059[129], stage058[132], stage057[137], stage056[149], stage055[188]}
   );
   gpc606_5 gpc606_5_1927(
      {stage055[68], stage055[69], stage055[70], stage055[71], stage055[72], stage055[73]},
      {stage057[12], stage057[13], stage057[14], stage057[15], stage057[16], stage057[17]},
      {stage059[130], stage058[133], stage057[138], stage056[150], stage055[189]}
   );
   gpc606_5 gpc606_5_1928(
      {stage055[74], stage055[75], stage055[76], stage055[77], stage055[78], stage055[79]},
      {stage057[18], stage057[19], stage057[20], stage057[21], stage057[22], stage057[23]},
      {stage059[131], stage058[134], stage057[139], stage056[151], stage055[190]}
   );
   gpc606_5 gpc606_5_1929(
      {stage055[80], stage055[81], stage055[82], stage055[83], stage055[84], stage055[85]},
      {stage057[24], stage057[25], stage057[26], stage057[27], stage057[28], stage057[29]},
      {stage059[132], stage058[135], stage057[140], stage056[152], stage055[191]}
   );
   gpc606_5 gpc606_5_1930(
      {stage055[86], stage055[87], stage055[88], stage055[89], stage055[90], stage055[91]},
      {stage057[30], stage057[31], stage057[32], stage057[33], stage057[34], stage057[35]},
      {stage059[133], stage058[136], stage057[141], stage056[153], stage055[192]}
   );
   gpc606_5 gpc606_5_1931(
      {stage055[92], stage055[93], stage055[94], stage055[95], stage055[96], stage055[97]},
      {stage057[36], stage057[37], stage057[38], stage057[39], stage057[40], stage057[41]},
      {stage059[134], stage058[137], stage057[142], stage056[154], stage055[193]}
   );
   gpc606_5 gpc606_5_1932(
      {stage055[98], stage055[99], stage055[100], stage055[101], stage055[102], stage055[103]},
      {stage057[42], stage057[43], stage057[44], stage057[45], stage057[46], stage057[47]},
      {stage059[135], stage058[138], stage057[143], stage056[155], stage055[194]}
   );
   gpc606_5 gpc606_5_1933(
      {stage055[104], stage055[105], stage055[106], stage055[107], stage055[108], stage055[109]},
      {stage057[48], stage057[49], stage057[50], stage057[51], stage057[52], stage057[53]},
      {stage059[136], stage058[139], stage057[144], stage056[156], stage055[195]}
   );
   gpc606_5 gpc606_5_1934(
      {stage055[110], stage055[111], stage055[112], stage055[113], stage055[114], stage055[115]},
      {stage057[54], stage057[55], stage057[56], stage057[57], stage057[58], stage057[59]},
      {stage059[137], stage058[140], stage057[145], stage056[157], stage055[196]}
   );
   gpc606_5 gpc606_5_1935(
      {stage055[116], stage055[117], stage055[118], stage055[119], stage055[120], stage055[121]},
      {stage057[60], stage057[61], stage057[62], stage057[63], stage057[64], stage057[65]},
      {stage059[138], stage058[141], stage057[146], stage056[158], stage055[197]}
   );
   gpc1406_5 gpc1406_5_1936(
      {stage055[122], stage055[123], stage055[124], stage055[125], stage055[126], stage055[127]},
      {stage057[66], stage057[67], stage057[68], stage057[69]},
      {stage058[0]},
      {stage059[139], stage058[142], stage057[147], stage056[159], stage055[198]}
   );
   gpc1_1 gpc1_1_1937(
      {stage056[18]},
      {stage056[160]}
   );
   gpc1_1 gpc1_1_1938(
      {stage056[19]},
      {stage056[161]}
   );
   gpc1_1 gpc1_1_1939(
      {stage056[20]},
      {stage056[162]}
   );
   gpc1_1 gpc1_1_1940(
      {stage056[21]},
      {stage056[163]}
   );
   gpc1_1 gpc1_1_1941(
      {stage056[22]},
      {stage056[164]}
   );
   gpc1_1 gpc1_1_1942(
      {stage056[23]},
      {stage056[165]}
   );
   gpc1_1 gpc1_1_1943(
      {stage056[24]},
      {stage056[166]}
   );
   gpc1_1 gpc1_1_1944(
      {stage056[25]},
      {stage056[167]}
   );
   gpc1_1 gpc1_1_1945(
      {stage056[26]},
      {stage056[168]}
   );
   gpc1_1 gpc1_1_1946(
      {stage056[27]},
      {stage056[169]}
   );
   gpc1_1 gpc1_1_1947(
      {stage056[28]},
      {stage056[170]}
   );
   gpc1_1 gpc1_1_1948(
      {stage056[29]},
      {stage056[171]}
   );
   gpc1_1 gpc1_1_1949(
      {stage056[30]},
      {stage056[172]}
   );
   gpc1_1 gpc1_1_1950(
      {stage056[31]},
      {stage056[173]}
   );
   gpc1_1 gpc1_1_1951(
      {stage056[32]},
      {stage056[174]}
   );
   gpc1_1 gpc1_1_1952(
      {stage056[33]},
      {stage056[175]}
   );
   gpc1_1 gpc1_1_1953(
      {stage056[34]},
      {stage056[176]}
   );
   gpc1_1 gpc1_1_1954(
      {stage056[35]},
      {stage056[177]}
   );
   gpc1_1 gpc1_1_1955(
      {stage056[36]},
      {stage056[178]}
   );
   gpc1_1 gpc1_1_1956(
      {stage056[37]},
      {stage056[179]}
   );
   gpc1_1 gpc1_1_1957(
      {stage056[38]},
      {stage056[180]}
   );
   gpc1_1 gpc1_1_1958(
      {stage056[39]},
      {stage056[181]}
   );
   gpc1_1 gpc1_1_1959(
      {stage056[40]},
      {stage056[182]}
   );
   gpc1_1 gpc1_1_1960(
      {stage056[41]},
      {stage056[183]}
   );
   gpc1_1 gpc1_1_1961(
      {stage056[42]},
      {stage056[184]}
   );
   gpc1_1 gpc1_1_1962(
      {stage056[43]},
      {stage056[185]}
   );
   gpc1_1 gpc1_1_1963(
      {stage056[44]},
      {stage056[186]}
   );
   gpc1_1 gpc1_1_1964(
      {stage056[45]},
      {stage056[187]}
   );
   gpc1_1 gpc1_1_1965(
      {stage056[46]},
      {stage056[188]}
   );
   gpc1_1 gpc1_1_1966(
      {stage056[47]},
      {stage056[189]}
   );
   gpc1_1 gpc1_1_1967(
      {stage056[48]},
      {stage056[190]}
   );
   gpc1_1 gpc1_1_1968(
      {stage056[49]},
      {stage056[191]}
   );
   gpc606_5 gpc606_5_1969(
      {stage056[50], stage056[51], stage056[52], stage056[53], stage056[54], stage056[55]},
      {stage058[1], stage058[2], stage058[3], stage058[4], stage058[5], stage058[6]},
      {stage060[128], stage059[140], stage058[143], stage057[148], stage056[192]}
   );
   gpc606_5 gpc606_5_1970(
      {stage056[56], stage056[57], stage056[58], stage056[59], stage056[60], stage056[61]},
      {stage058[7], stage058[8], stage058[9], stage058[10], stage058[11], stage058[12]},
      {stage060[129], stage059[141], stage058[144], stage057[149], stage056[193]}
   );
   gpc606_5 gpc606_5_1971(
      {stage056[62], stage056[63], stage056[64], stage056[65], stage056[66], stage056[67]},
      {stage058[13], stage058[14], stage058[15], stage058[16], stage058[17], stage058[18]},
      {stage060[130], stage059[142], stage058[145], stage057[150], stage056[194]}
   );
   gpc606_5 gpc606_5_1972(
      {stage056[68], stage056[69], stage056[70], stage056[71], stage056[72], stage056[73]},
      {stage058[19], stage058[20], stage058[21], stage058[22], stage058[23], stage058[24]},
      {stage060[131], stage059[143], stage058[146], stage057[151], stage056[195]}
   );
   gpc606_5 gpc606_5_1973(
      {stage056[74], stage056[75], stage056[76], stage056[77], stage056[78], stage056[79]},
      {stage058[25], stage058[26], stage058[27], stage058[28], stage058[29], stage058[30]},
      {stage060[132], stage059[144], stage058[147], stage057[152], stage056[196]}
   );
   gpc606_5 gpc606_5_1974(
      {stage056[80], stage056[81], stage056[82], stage056[83], stage056[84], stage056[85]},
      {stage058[31], stage058[32], stage058[33], stage058[34], stage058[35], stage058[36]},
      {stage060[133], stage059[145], stage058[148], stage057[153], stage056[197]}
   );
   gpc606_5 gpc606_5_1975(
      {stage056[86], stage056[87], stage056[88], stage056[89], stage056[90], stage056[91]},
      {stage058[37], stage058[38], stage058[39], stage058[40], stage058[41], stage058[42]},
      {stage060[134], stage059[146], stage058[149], stage057[154], stage056[198]}
   );
   gpc606_5 gpc606_5_1976(
      {stage056[92], stage056[93], stage056[94], stage056[95], stage056[96], stage056[97]},
      {stage058[43], stage058[44], stage058[45], stage058[46], stage058[47], stage058[48]},
      {stage060[135], stage059[147], stage058[150], stage057[155], stage056[199]}
   );
   gpc606_5 gpc606_5_1977(
      {stage056[98], stage056[99], stage056[100], stage056[101], stage056[102], stage056[103]},
      {stage058[49], stage058[50], stage058[51], stage058[52], stage058[53], stage058[54]},
      {stage060[136], stage059[148], stage058[151], stage057[156], stage056[200]}
   );
   gpc606_5 gpc606_5_1978(
      {stage056[104], stage056[105], stage056[106], stage056[107], stage056[108], stage056[109]},
      {stage058[55], stage058[56], stage058[57], stage058[58], stage058[59], stage058[60]},
      {stage060[137], stage059[149], stage058[152], stage057[157], stage056[201]}
   );
   gpc606_5 gpc606_5_1979(
      {stage056[110], stage056[111], stage056[112], stage056[113], stage056[114], stage056[115]},
      {stage058[61], stage058[62], stage058[63], stage058[64], stage058[65], stage058[66]},
      {stage060[138], stage059[150], stage058[153], stage057[158], stage056[202]}
   );
   gpc606_5 gpc606_5_1980(
      {stage056[116], stage056[117], stage056[118], stage056[119], stage056[120], stage056[121]},
      {stage058[67], stage058[68], stage058[69], stage058[70], stage058[71], stage058[72]},
      {stage060[139], stage059[151], stage058[154], stage057[159], stage056[203]}
   );
   gpc606_5 gpc606_5_1981(
      {stage056[122], stage056[123], stage056[124], stage056[125], stage056[126], stage056[127]},
      {stage058[73], stage058[74], stage058[75], stage058[76], stage058[77], stage058[78]},
      {stage060[140], stage059[152], stage058[155], stage057[160], stage056[204]}
   );
   gpc1_1 gpc1_1_1982(
      {stage057[70]},
      {stage057[161]}
   );
   gpc1_1 gpc1_1_1983(
      {stage057[71]},
      {stage057[162]}
   );
   gpc1_1 gpc1_1_1984(
      {stage057[72]},
      {stage057[163]}
   );
   gpc1_1 gpc1_1_1985(
      {stage057[73]},
      {stage057[164]}
   );
   gpc1_1 gpc1_1_1986(
      {stage057[74]},
      {stage057[165]}
   );
   gpc1_1 gpc1_1_1987(
      {stage057[75]},
      {stage057[166]}
   );
   gpc1_1 gpc1_1_1988(
      {stage057[76]},
      {stage057[167]}
   );
   gpc1_1 gpc1_1_1989(
      {stage057[77]},
      {stage057[168]}
   );
   gpc1_1 gpc1_1_1990(
      {stage057[78]},
      {stage057[169]}
   );
   gpc1_1 gpc1_1_1991(
      {stage057[79]},
      {stage057[170]}
   );
   gpc1_1 gpc1_1_1992(
      {stage057[80]},
      {stage057[171]}
   );
   gpc1_1 gpc1_1_1993(
      {stage057[81]},
      {stage057[172]}
   );
   gpc1_1 gpc1_1_1994(
      {stage057[82]},
      {stage057[173]}
   );
   gpc1_1 gpc1_1_1995(
      {stage057[83]},
      {stage057[174]}
   );
   gpc1_1 gpc1_1_1996(
      {stage057[84]},
      {stage057[175]}
   );
   gpc1_1 gpc1_1_1997(
      {stage057[85]},
      {stage057[176]}
   );
   gpc606_5 gpc606_5_1998(
      {stage057[86], stage057[87], stage057[88], stage057[89], stage057[90], stage057[91]},
      {stage059[0], stage059[1], stage059[2], stage059[3], stage059[4], stage059[5]},
      {stage061[128], stage060[141], stage059[153], stage058[156], stage057[177]}
   );
   gpc606_5 gpc606_5_1999(
      {stage057[92], stage057[93], stage057[94], stage057[95], stage057[96], stage057[97]},
      {stage059[6], stage059[7], stage059[8], stage059[9], stage059[10], stage059[11]},
      {stage061[129], stage060[142], stage059[154], stage058[157], stage057[178]}
   );
   gpc606_5 gpc606_5_2000(
      {stage057[98], stage057[99], stage057[100], stage057[101], stage057[102], stage057[103]},
      {stage059[12], stage059[13], stage059[14], stage059[15], stage059[16], stage059[17]},
      {stage061[130], stage060[143], stage059[155], stage058[158], stage057[179]}
   );
   gpc606_5 gpc606_5_2001(
      {stage057[104], stage057[105], stage057[106], stage057[107], stage057[108], stage057[109]},
      {stage059[18], stage059[19], stage059[20], stage059[21], stage059[22], stage059[23]},
      {stage061[131], stage060[144], stage059[156], stage058[159], stage057[180]}
   );
   gpc606_5 gpc606_5_2002(
      {stage057[110], stage057[111], stage057[112], stage057[113], stage057[114], stage057[115]},
      {stage059[24], stage059[25], stage059[26], stage059[27], stage059[28], stage059[29]},
      {stage061[132], stage060[145], stage059[157], stage058[160], stage057[181]}
   );
   gpc606_5 gpc606_5_2003(
      {stage057[116], stage057[117], stage057[118], stage057[119], stage057[120], stage057[121]},
      {stage059[30], stage059[31], stage059[32], stage059[33], stage059[34], stage059[35]},
      {stage061[133], stage060[146], stage059[158], stage058[161], stage057[182]}
   );
   gpc606_5 gpc606_5_2004(
      {stage057[122], stage057[123], stage057[124], stage057[125], stage057[126], stage057[127]},
      {stage059[36], stage059[37], stage059[38], stage059[39], stage059[40], stage059[41]},
      {stage061[134], stage060[147], stage059[159], stage058[162], stage057[183]}
   );
   gpc1_1 gpc1_1_2005(
      {stage058[79]},
      {stage058[163]}
   );
   gpc1_1 gpc1_1_2006(
      {stage058[80]},
      {stage058[164]}
   );
   gpc1_1 gpc1_1_2007(
      {stage058[81]},
      {stage058[165]}
   );
   gpc1_1 gpc1_1_2008(
      {stage058[82]},
      {stage058[166]}
   );
   gpc1_1 gpc1_1_2009(
      {stage058[83]},
      {stage058[167]}
   );
   gpc1_1 gpc1_1_2010(
      {stage058[84]},
      {stage058[168]}
   );
   gpc1_1 gpc1_1_2011(
      {stage058[85]},
      {stage058[169]}
   );
   gpc1_1 gpc1_1_2012(
      {stage058[86]},
      {stage058[170]}
   );
   gpc1_1 gpc1_1_2013(
      {stage058[87]},
      {stage058[171]}
   );
   gpc615_5 gpc615_5_2014(
      {stage058[88], stage058[89], stage058[90], stage058[91], stage058[92]},
      {stage059[42]},
      {stage060[0], stage060[1], stage060[2], stage060[3], stage060[4], stage060[5]},
      {stage062[128], stage061[135], stage060[148], stage059[160], stage058[172]}
   );
   gpc615_5 gpc615_5_2015(
      {stage058[93], stage058[94], stage058[95], stage058[96], stage058[97]},
      {stage059[43]},
      {stage060[6], stage060[7], stage060[8], stage060[9], stage060[10], stage060[11]},
      {stage062[129], stage061[136], stage060[149], stage059[161], stage058[173]}
   );
   gpc615_5 gpc615_5_2016(
      {stage058[98], stage058[99], stage058[100], stage058[101], stage058[102]},
      {stage059[44]},
      {stage060[12], stage060[13], stage060[14], stage060[15], stage060[16], stage060[17]},
      {stage062[130], stage061[137], stage060[150], stage059[162], stage058[174]}
   );
   gpc615_5 gpc615_5_2017(
      {stage058[103], stage058[104], stage058[105], stage058[106], stage058[107]},
      {stage059[45]},
      {stage060[18], stage060[19], stage060[20], stage060[21], stage060[22], stage060[23]},
      {stage062[131], stage061[138], stage060[151], stage059[163], stage058[175]}
   );
   gpc615_5 gpc615_5_2018(
      {stage058[108], stage058[109], stage058[110], stage058[111], stage058[112]},
      {stage059[46]},
      {stage060[24], stage060[25], stage060[26], stage060[27], stage060[28], stage060[29]},
      {stage062[132], stage061[139], stage060[152], stage059[164], stage058[176]}
   );
   gpc615_5 gpc615_5_2019(
      {stage058[113], stage058[114], stage058[115], stage058[116], stage058[117]},
      {stage059[47]},
      {stage060[30], stage060[31], stage060[32], stage060[33], stage060[34], stage060[35]},
      {stage062[133], stage061[140], stage060[153], stage059[165], stage058[177]}
   );
   gpc615_5 gpc615_5_2020(
      {stage058[118], stage058[119], stage058[120], stage058[121], stage058[122]},
      {stage059[48]},
      {stage060[36], stage060[37], stage060[38], stage060[39], stage060[40], stage060[41]},
      {stage062[134], stage061[141], stage060[154], stage059[166], stage058[178]}
   );
   gpc615_5 gpc615_5_2021(
      {stage058[123], stage058[124], stage058[125], stage058[126], stage058[127]},
      {stage059[49]},
      {stage060[42], stage060[43], stage060[44], stage060[45], stage060[46], stage060[47]},
      {stage062[135], stage061[142], stage060[155], stage059[167], stage058[179]}
   );
   gpc1_1 gpc1_1_2022(
      {stage059[50]},
      {stage059[168]}
   );
   gpc1_1 gpc1_1_2023(
      {stage059[51]},
      {stage059[169]}
   );
   gpc1_1 gpc1_1_2024(
      {stage059[52]},
      {stage059[170]}
   );
   gpc1_1 gpc1_1_2025(
      {stage059[53]},
      {stage059[171]}
   );
   gpc1_1 gpc1_1_2026(
      {stage059[54]},
      {stage059[172]}
   );
   gpc1_1 gpc1_1_2027(
      {stage059[55]},
      {stage059[173]}
   );
   gpc1_1 gpc1_1_2028(
      {stage059[56]},
      {stage059[174]}
   );
   gpc1_1 gpc1_1_2029(
      {stage059[57]},
      {stage059[175]}
   );
   gpc1_1 gpc1_1_2030(
      {stage059[58]},
      {stage059[176]}
   );
   gpc1_1 gpc1_1_2031(
      {stage059[59]},
      {stage059[177]}
   );
   gpc1_1 gpc1_1_2032(
      {stage059[60]},
      {stage059[178]}
   );
   gpc1_1 gpc1_1_2033(
      {stage059[61]},
      {stage059[179]}
   );
   gpc1_1 gpc1_1_2034(
      {stage059[62]},
      {stage059[180]}
   );
   gpc1_1 gpc1_1_2035(
      {stage059[63]},
      {stage059[181]}
   );
   gpc1_1 gpc1_1_2036(
      {stage059[64]},
      {stage059[182]}
   );
   gpc1_1 gpc1_1_2037(
      {stage059[65]},
      {stage059[183]}
   );
   gpc1_1 gpc1_1_2038(
      {stage059[66]},
      {stage059[184]}
   );
   gpc1_1 gpc1_1_2039(
      {stage059[67]},
      {stage059[185]}
   );
   gpc1_1 gpc1_1_2040(
      {stage059[68]},
      {stage059[186]}
   );
   gpc1_1 gpc1_1_2041(
      {stage059[69]},
      {stage059[187]}
   );
   gpc1_1 gpc1_1_2042(
      {stage059[70]},
      {stage059[188]}
   );
   gpc1_1 gpc1_1_2043(
      {stage059[71]},
      {stage059[189]}
   );
   gpc1_1 gpc1_1_2044(
      {stage059[72]},
      {stage059[190]}
   );
   gpc1_1 gpc1_1_2045(
      {stage059[73]},
      {stage059[191]}
   );
   gpc1_1 gpc1_1_2046(
      {stage059[74]},
      {stage059[192]}
   );
   gpc1_1 gpc1_1_2047(
      {stage059[75]},
      {stage059[193]}
   );
   gpc1_1 gpc1_1_2048(
      {stage059[76]},
      {stage059[194]}
   );
   gpc1_1 gpc1_1_2049(
      {stage059[77]},
      {stage059[195]}
   );
   gpc1_1 gpc1_1_2050(
      {stage059[78]},
      {stage059[196]}
   );
   gpc1_1 gpc1_1_2051(
      {stage059[79]},
      {stage059[197]}
   );
   gpc1_1 gpc1_1_2052(
      {stage059[80]},
      {stage059[198]}
   );
   gpc1_1 gpc1_1_2053(
      {stage059[81]},
      {stage059[199]}
   );
   gpc1_1 gpc1_1_2054(
      {stage059[82]},
      {stage059[200]}
   );
   gpc1_1 gpc1_1_2055(
      {stage059[83]},
      {stage059[201]}
   );
   gpc1_1 gpc1_1_2056(
      {stage059[84]},
      {stage059[202]}
   );
   gpc1_1 gpc1_1_2057(
      {stage059[85]},
      {stage059[203]}
   );
   gpc1_1 gpc1_1_2058(
      {stage059[86]},
      {stage059[204]}
   );
   gpc1_1 gpc1_1_2059(
      {stage059[87]},
      {stage059[205]}
   );
   gpc1_1 gpc1_1_2060(
      {stage059[88]},
      {stage059[206]}
   );
   gpc1_1 gpc1_1_2061(
      {stage059[89]},
      {stage059[207]}
   );
   gpc1_1 gpc1_1_2062(
      {stage059[90]},
      {stage059[208]}
   );
   gpc1_1 gpc1_1_2063(
      {stage059[91]},
      {stage059[209]}
   );
   gpc606_5 gpc606_5_2064(
      {stage059[92], stage059[93], stage059[94], stage059[95], stage059[96], stage059[97]},
      {stage061[0], stage061[1], stage061[2], stage061[3], stage061[4], stage061[5]},
      {stage063[128], stage062[136], stage061[143], stage060[156], stage059[210]}
   );
   gpc606_5 gpc606_5_2065(
      {stage059[98], stage059[99], stage059[100], stage059[101], stage059[102], stage059[103]},
      {stage061[6], stage061[7], stage061[8], stage061[9], stage061[10], stage061[11]},
      {stage063[129], stage062[137], stage061[144], stage060[157], stage059[211]}
   );
   gpc606_5 gpc606_5_2066(
      {stage059[104], stage059[105], stage059[106], stage059[107], stage059[108], stage059[109]},
      {stage061[12], stage061[13], stage061[14], stage061[15], stage061[16], stage061[17]},
      {stage063[130], stage062[138], stage061[145], stage060[158], stage059[212]}
   );
   gpc606_5 gpc606_5_2067(
      {stage059[110], stage059[111], stage059[112], stage059[113], stage059[114], stage059[115]},
      {stage061[18], stage061[19], stage061[20], stage061[21], stage061[22], stage061[23]},
      {stage063[131], stage062[139], stage061[146], stage060[159], stage059[213]}
   );
   gpc606_5 gpc606_5_2068(
      {stage059[116], stage059[117], stage059[118], stage059[119], stage059[120], stage059[121]},
      {stage061[24], stage061[25], stage061[26], stage061[27], stage061[28], stage061[29]},
      {stage063[132], stage062[140], stage061[147], stage060[160], stage059[214]}
   );
   gpc606_5 gpc606_5_2069(
      {stage059[122], stage059[123], stage059[124], stage059[125], stage059[126], stage059[127]},
      {stage061[30], stage061[31], stage061[32], stage061[33], stage061[34], stage061[35]},
      {stage063[133], stage062[141], stage061[148], stage060[161], stage059[215]}
   );
   gpc1_1 gpc1_1_2070(
      {stage060[48]},
      {stage060[162]}
   );
   gpc1_1 gpc1_1_2071(
      {stage060[49]},
      {stage060[163]}
   );
   gpc1_1 gpc1_1_2072(
      {stage060[50]},
      {stage060[164]}
   );
   gpc1_1 gpc1_1_2073(
      {stage060[51]},
      {stage060[165]}
   );
   gpc1_1 gpc1_1_2074(
      {stage060[52]},
      {stage060[166]}
   );
   gpc1_1 gpc1_1_2075(
      {stage060[53]},
      {stage060[167]}
   );
   gpc1_1 gpc1_1_2076(
      {stage060[54]},
      {stage060[168]}
   );
   gpc1_1 gpc1_1_2077(
      {stage060[55]},
      {stage060[169]}
   );
   gpc1_1 gpc1_1_2078(
      {stage060[56]},
      {stage060[170]}
   );
   gpc1_1 gpc1_1_2079(
      {stage060[57]},
      {stage060[171]}
   );
   gpc1_1 gpc1_1_2080(
      {stage060[58]},
      {stage060[172]}
   );
   gpc1_1 gpc1_1_2081(
      {stage060[59]},
      {stage060[173]}
   );
   gpc1_1 gpc1_1_2082(
      {stage060[60]},
      {stage060[174]}
   );
   gpc1_1 gpc1_1_2083(
      {stage060[61]},
      {stage060[175]}
   );
   gpc1_1 gpc1_1_2084(
      {stage060[62]},
      {stage060[176]}
   );
   gpc615_5 gpc615_5_2085(
      {stage060[63], stage060[64], stage060[65], stage060[66], stage060[67]},
      {stage061[36]},
      {stage062[0], stage062[1], stage062[2], stage062[3], stage062[4], stage062[5]},
      {stage064[128], stage063[134], stage062[142], stage061[149], stage060[177]}
   );
   gpc615_5 gpc615_5_2086(
      {stage060[68], stage060[69], stage060[70], stage060[71], stage060[72]},
      {stage061[37]},
      {stage062[6], stage062[7], stage062[8], stage062[9], stage062[10], stage062[11]},
      {stage064[129], stage063[135], stage062[143], stage061[150], stage060[178]}
   );
   gpc615_5 gpc615_5_2087(
      {stage060[73], stage060[74], stage060[75], stage060[76], stage060[77]},
      {stage061[38]},
      {stage062[12], stage062[13], stage062[14], stage062[15], stage062[16], stage062[17]},
      {stage064[130], stage063[136], stage062[144], stage061[151], stage060[179]}
   );
   gpc615_5 gpc615_5_2088(
      {stage060[78], stage060[79], stage060[80], stage060[81], stage060[82]},
      {stage061[39]},
      {stage062[18], stage062[19], stage062[20], stage062[21], stage062[22], stage062[23]},
      {stage064[131], stage063[137], stage062[145], stage061[152], stage060[180]}
   );
   gpc615_5 gpc615_5_2089(
      {stage060[83], stage060[84], stage060[85], stage060[86], stage060[87]},
      {stage061[40]},
      {stage062[24], stage062[25], stage062[26], stage062[27], stage062[28], stage062[29]},
      {stage064[132], stage063[138], stage062[146], stage061[153], stage060[181]}
   );
   gpc615_5 gpc615_5_2090(
      {stage060[88], stage060[89], stage060[90], stage060[91], stage060[92]},
      {stage061[41]},
      {stage062[30], stage062[31], stage062[32], stage062[33], stage062[34], stage062[35]},
      {stage064[133], stage063[139], stage062[147], stage061[154], stage060[182]}
   );
   gpc615_5 gpc615_5_2091(
      {stage060[93], stage060[94], stage060[95], stage060[96], stage060[97]},
      {stage061[42]},
      {stage062[36], stage062[37], stage062[38], stage062[39], stage062[40], stage062[41]},
      {stage064[134], stage063[140], stage062[148], stage061[155], stage060[183]}
   );
   gpc615_5 gpc615_5_2092(
      {stage060[98], stage060[99], stage060[100], stage060[101], stage060[102]},
      {stage061[43]},
      {stage062[42], stage062[43], stage062[44], stage062[45], stage062[46], stage062[47]},
      {stage064[135], stage063[141], stage062[149], stage061[156], stage060[184]}
   );
   gpc615_5 gpc615_5_2093(
      {stage060[103], stage060[104], stage060[105], stage060[106], stage060[107]},
      {stage061[44]},
      {stage062[48], stage062[49], stage062[50], stage062[51], stage062[52], stage062[53]},
      {stage064[136], stage063[142], stage062[150], stage061[157], stage060[185]}
   );
   gpc615_5 gpc615_5_2094(
      {stage060[108], stage060[109], stage060[110], stage060[111], stage060[112]},
      {stage061[45]},
      {stage062[54], stage062[55], stage062[56], stage062[57], stage062[58], stage062[59]},
      {stage064[137], stage063[143], stage062[151], stage061[158], stage060[186]}
   );
   gpc615_5 gpc615_5_2095(
      {stage060[113], stage060[114], stage060[115], stage060[116], stage060[117]},
      {stage061[46]},
      {stage062[60], stage062[61], stage062[62], stage062[63], stage062[64], stage062[65]},
      {stage064[138], stage063[144], stage062[152], stage061[159], stage060[187]}
   );
   gpc615_5 gpc615_5_2096(
      {stage060[118], stage060[119], stage060[120], stage060[121], stage060[122]},
      {stage061[47]},
      {stage062[66], stage062[67], stage062[68], stage062[69], stage062[70], stage062[71]},
      {stage064[139], stage063[145], stage062[153], stage061[160], stage060[188]}
   );
   gpc615_5 gpc615_5_2097(
      {stage060[123], stage060[124], stage060[125], stage060[126], stage060[127]},
      {stage061[48]},
      {stage062[72], stage062[73], stage062[74], stage062[75], stage062[76], stage062[77]},
      {stage064[140], stage063[146], stage062[154], stage061[161], stage060[189]}
   );
   gpc1_1 gpc1_1_2098(
      {stage061[49]},
      {stage061[162]}
   );
   gpc1_1 gpc1_1_2099(
      {stage061[50]},
      {stage061[163]}
   );
   gpc1_1 gpc1_1_2100(
      {stage061[51]},
      {stage061[164]}
   );
   gpc1_1 gpc1_1_2101(
      {stage061[52]},
      {stage061[165]}
   );
   gpc1_1 gpc1_1_2102(
      {stage061[53]},
      {stage061[166]}
   );
   gpc1_1 gpc1_1_2103(
      {stage061[54]},
      {stage061[167]}
   );
   gpc1_1 gpc1_1_2104(
      {stage061[55]},
      {stage061[168]}
   );
   gpc1_1 gpc1_1_2105(
      {stage061[56]},
      {stage061[169]}
   );
   gpc1_1 gpc1_1_2106(
      {stage061[57]},
      {stage061[170]}
   );
   gpc1_1 gpc1_1_2107(
      {stage061[58]},
      {stage061[171]}
   );
   gpc1_1 gpc1_1_2108(
      {stage061[59]},
      {stage061[172]}
   );
   gpc1_1 gpc1_1_2109(
      {stage061[60]},
      {stage061[173]}
   );
   gpc1_1 gpc1_1_2110(
      {stage061[61]},
      {stage061[174]}
   );
   gpc1_1 gpc1_1_2111(
      {stage061[62]},
      {stage061[175]}
   );
   gpc615_5 gpc615_5_2112(
      {stage061[63], stage061[64], stage061[65], stage061[66], stage061[67]},
      {stage062[78]},
      {stage063[0], stage063[1], stage063[2], stage063[3], stage063[4], stage063[5]},
      {stage065[128], stage064[141], stage063[147], stage062[155], stage061[176]}
   );
   gpc615_5 gpc615_5_2113(
      {stage061[68], stage061[69], stage061[70], stage061[71], stage061[72]},
      {stage062[79]},
      {stage063[6], stage063[7], stage063[8], stage063[9], stage063[10], stage063[11]},
      {stage065[129], stage064[142], stage063[148], stage062[156], stage061[177]}
   );
   gpc615_5 gpc615_5_2114(
      {stage061[73], stage061[74], stage061[75], stage061[76], stage061[77]},
      {stage062[80]},
      {stage063[12], stage063[13], stage063[14], stage063[15], stage063[16], stage063[17]},
      {stage065[130], stage064[143], stage063[149], stage062[157], stage061[178]}
   );
   gpc615_5 gpc615_5_2115(
      {stage061[78], stage061[79], stage061[80], stage061[81], stage061[82]},
      {stage062[81]},
      {stage063[18], stage063[19], stage063[20], stage063[21], stage063[22], stage063[23]},
      {stage065[131], stage064[144], stage063[150], stage062[158], stage061[179]}
   );
   gpc615_5 gpc615_5_2116(
      {stage061[83], stage061[84], stage061[85], stage061[86], stage061[87]},
      {stage062[82]},
      {stage063[24], stage063[25], stage063[26], stage063[27], stage063[28], stage063[29]},
      {stage065[132], stage064[145], stage063[151], stage062[159], stage061[180]}
   );
   gpc615_5 gpc615_5_2117(
      {stage061[88], stage061[89], stage061[90], stage061[91], stage061[92]},
      {stage062[83]},
      {stage063[30], stage063[31], stage063[32], stage063[33], stage063[34], stage063[35]},
      {stage065[133], stage064[146], stage063[152], stage062[160], stage061[181]}
   );
   gpc615_5 gpc615_5_2118(
      {stage061[93], stage061[94], stage061[95], stage061[96], stage061[97]},
      {stage062[84]},
      {stage063[36], stage063[37], stage063[38], stage063[39], stage063[40], stage063[41]},
      {stage065[134], stage064[147], stage063[153], stage062[161], stage061[182]}
   );
   gpc615_5 gpc615_5_2119(
      {stage061[98], stage061[99], stage061[100], stage061[101], stage061[102]},
      {stage062[85]},
      {stage063[42], stage063[43], stage063[44], stage063[45], stage063[46], stage063[47]},
      {stage065[135], stage064[148], stage063[154], stage062[162], stage061[183]}
   );
   gpc615_5 gpc615_5_2120(
      {stage061[103], stage061[104], stage061[105], stage061[106], stage061[107]},
      {stage062[86]},
      {stage063[48], stage063[49], stage063[50], stage063[51], stage063[52], stage063[53]},
      {stage065[136], stage064[149], stage063[155], stage062[163], stage061[184]}
   );
   gpc615_5 gpc615_5_2121(
      {stage061[108], stage061[109], stage061[110], stage061[111], stage061[112]},
      {stage062[87]},
      {stage063[54], stage063[55], stage063[56], stage063[57], stage063[58], stage063[59]},
      {stage065[137], stage064[150], stage063[156], stage062[164], stage061[185]}
   );
   gpc615_5 gpc615_5_2122(
      {stage061[113], stage061[114], stage061[115], stage061[116], stage061[117]},
      {stage062[88]},
      {stage063[60], stage063[61], stage063[62], stage063[63], stage063[64], stage063[65]},
      {stage065[138], stage064[151], stage063[157], stage062[165], stage061[186]}
   );
   gpc615_5 gpc615_5_2123(
      {stage061[118], stage061[119], stage061[120], stage061[121], stage061[122]},
      {stage062[89]},
      {stage063[66], stage063[67], stage063[68], stage063[69], stage063[70], stage063[71]},
      {stage065[139], stage064[152], stage063[158], stage062[166], stage061[187]}
   );
   gpc615_5 gpc615_5_2124(
      {stage061[123], stage061[124], stage061[125], stage061[126], stage061[127]},
      {stage062[90]},
      {stage063[72], stage063[73], stage063[74], stage063[75], stage063[76], stage063[77]},
      {stage065[140], stage064[153], stage063[159], stage062[167], stage061[188]}
   );
   gpc1_1 gpc1_1_2125(
      {stage062[91]},
      {stage062[168]}
   );
   gpc1_1 gpc1_1_2126(
      {stage062[92]},
      {stage062[169]}
   );
   gpc1_1 gpc1_1_2127(
      {stage062[93]},
      {stage062[170]}
   );
   gpc1_1 gpc1_1_2128(
      {stage062[94]},
      {stage062[171]}
   );
   gpc1_1 gpc1_1_2129(
      {stage062[95]},
      {stage062[172]}
   );
   gpc1_1 gpc1_1_2130(
      {stage062[96]},
      {stage062[173]}
   );
   gpc1_1 gpc1_1_2131(
      {stage062[97]},
      {stage062[174]}
   );
   gpc1_1 gpc1_1_2132(
      {stage062[98]},
      {stage062[175]}
   );
   gpc1_1 gpc1_1_2133(
      {stage062[99]},
      {stage062[176]}
   );
   gpc1_1 gpc1_1_2134(
      {stage062[100]},
      {stage062[177]}
   );
   gpc1_1 gpc1_1_2135(
      {stage062[101]},
      {stage062[178]}
   );
   gpc1_1 gpc1_1_2136(
      {stage062[102]},
      {stage062[179]}
   );
   gpc1_1 gpc1_1_2137(
      {stage062[103]},
      {stage062[180]}
   );
   gpc1_1 gpc1_1_2138(
      {stage062[104]},
      {stage062[181]}
   );
   gpc1_1 gpc1_1_2139(
      {stage062[105]},
      {stage062[182]}
   );
   gpc1_1 gpc1_1_2140(
      {stage062[106]},
      {stage062[183]}
   );
   gpc1_1 gpc1_1_2141(
      {stage062[107]},
      {stage062[184]}
   );
   gpc615_5 gpc615_5_2142(
      {stage062[108], stage062[109], stage062[110], stage062[111], stage062[112]},
      {stage063[78]},
      {stage064[0], stage064[1], stage064[2], stage064[3], stage064[4], stage064[5]},
      {stage066[128], stage065[141], stage064[154], stage063[160], stage062[185]}
   );
   gpc615_5 gpc615_5_2143(
      {stage062[113], stage062[114], stage062[115], stage062[116], stage062[117]},
      {stage063[79]},
      {stage064[6], stage064[7], stage064[8], stage064[9], stage064[10], stage064[11]},
      {stage066[129], stage065[142], stage064[155], stage063[161], stage062[186]}
   );
   gpc615_5 gpc615_5_2144(
      {stage062[118], stage062[119], stage062[120], stage062[121], stage062[122]},
      {stage063[80]},
      {stage064[12], stage064[13], stage064[14], stage064[15], stage064[16], stage064[17]},
      {stage066[130], stage065[143], stage064[156], stage063[162], stage062[187]}
   );
   gpc615_5 gpc615_5_2145(
      {stage062[123], stage062[124], stage062[125], stage062[126], stage062[127]},
      {stage063[81]},
      {stage064[18], stage064[19], stage064[20], stage064[21], stage064[22], stage064[23]},
      {stage066[131], stage065[144], stage064[157], stage063[163], stage062[188]}
   );
   gpc1_1 gpc1_1_2146(
      {stage063[82]},
      {stage063[164]}
   );
   gpc1_1 gpc1_1_2147(
      {stage063[83]},
      {stage063[165]}
   );
   gpc1_1 gpc1_1_2148(
      {stage063[84]},
      {stage063[166]}
   );
   gpc1_1 gpc1_1_2149(
      {stage063[85]},
      {stage063[167]}
   );
   gpc606_5 gpc606_5_2150(
      {stage063[86], stage063[87], stage063[88], stage063[89], stage063[90], stage063[91]},
      {stage065[0], stage065[1], stage065[2], stage065[3], stage065[4], stage065[5]},
      {stage067[128], stage066[132], stage065[145], stage064[158], stage063[168]}
   );
   gpc606_5 gpc606_5_2151(
      {stage063[92], stage063[93], stage063[94], stage063[95], stage063[96], stage063[97]},
      {stage065[6], stage065[7], stage065[8], stage065[9], stage065[10], stage065[11]},
      {stage067[129], stage066[133], stage065[146], stage064[159], stage063[169]}
   );
   gpc606_5 gpc606_5_2152(
      {stage063[98], stage063[99], stage063[100], stage063[101], stage063[102], stage063[103]},
      {stage065[12], stage065[13], stage065[14], stage065[15], stage065[16], stage065[17]},
      {stage067[130], stage066[134], stage065[147], stage064[160], stage063[170]}
   );
   gpc606_5 gpc606_5_2153(
      {stage063[104], stage063[105], stage063[106], stage063[107], stage063[108], stage063[109]},
      {stage065[18], stage065[19], stage065[20], stage065[21], stage065[22], stage065[23]},
      {stage067[131], stage066[135], stage065[148], stage064[161], stage063[171]}
   );
   gpc606_5 gpc606_5_2154(
      {stage063[110], stage063[111], stage063[112], stage063[113], stage063[114], stage063[115]},
      {stage065[24], stage065[25], stage065[26], stage065[27], stage065[28], stage065[29]},
      {stage067[132], stage066[136], stage065[149], stage064[162], stage063[172]}
   );
   gpc606_5 gpc606_5_2155(
      {stage063[116], stage063[117], stage063[118], stage063[119], stage063[120], stage063[121]},
      {stage065[30], stage065[31], stage065[32], stage065[33], stage065[34], stage065[35]},
      {stage067[133], stage066[137], stage065[150], stage064[163], stage063[173]}
   );
   gpc606_5 gpc606_5_2156(
      {stage063[122], stage063[123], stage063[124], stage063[125], stage063[126], stage063[127]},
      {stage065[36], stage065[37], stage065[38], stage065[39], stage065[40], stage065[41]},
      {stage067[134], stage066[138], stage065[151], stage064[164], stage063[174]}
   );
   gpc1_1 gpc1_1_2157(
      {stage064[24]},
      {stage064[165]}
   );
   gpc1_1 gpc1_1_2158(
      {stage064[25]},
      {stage064[166]}
   );
   gpc1_1 gpc1_1_2159(
      {stage064[26]},
      {stage064[167]}
   );
   gpc1_1 gpc1_1_2160(
      {stage064[27]},
      {stage064[168]}
   );
   gpc1_1 gpc1_1_2161(
      {stage064[28]},
      {stage064[169]}
   );
   gpc1_1 gpc1_1_2162(
      {stage064[29]},
      {stage064[170]}
   );
   gpc1_1 gpc1_1_2163(
      {stage064[30]},
      {stage064[171]}
   );
   gpc1_1 gpc1_1_2164(
      {stage064[31]},
      {stage064[172]}
   );
   gpc1_1 gpc1_1_2165(
      {stage064[32]},
      {stage064[173]}
   );
   gpc1_1 gpc1_1_2166(
      {stage064[33]},
      {stage064[174]}
   );
   gpc1_1 gpc1_1_2167(
      {stage064[34]},
      {stage064[175]}
   );
   gpc1_1 gpc1_1_2168(
      {stage064[35]},
      {stage064[176]}
   );
   gpc1_1 gpc1_1_2169(
      {stage064[36]},
      {stage064[177]}
   );
   gpc1_1 gpc1_1_2170(
      {stage064[37]},
      {stage064[178]}
   );
   gpc1_1 gpc1_1_2171(
      {stage064[38]},
      {stage064[179]}
   );
   gpc1_1 gpc1_1_2172(
      {stage064[39]},
      {stage064[180]}
   );
   gpc1_1 gpc1_1_2173(
      {stage064[40]},
      {stage064[181]}
   );
   gpc1_1 gpc1_1_2174(
      {stage064[41]},
      {stage064[182]}
   );
   gpc1_1 gpc1_1_2175(
      {stage064[42]},
      {stage064[183]}
   );
   gpc1_1 gpc1_1_2176(
      {stage064[43]},
      {stage064[184]}
   );
   gpc1_1 gpc1_1_2177(
      {stage064[44]},
      {stage064[185]}
   );
   gpc1_1 gpc1_1_2178(
      {stage064[45]},
      {stage064[186]}
   );
   gpc1_1 gpc1_1_2179(
      {stage064[46]},
      {stage064[187]}
   );
   gpc1_1 gpc1_1_2180(
      {stage064[47]},
      {stage064[188]}
   );
   gpc1_1 gpc1_1_2181(
      {stage064[48]},
      {stage064[189]}
   );
   gpc1_1 gpc1_1_2182(
      {stage064[49]},
      {stage064[190]}
   );
   gpc1_1 gpc1_1_2183(
      {stage064[50]},
      {stage064[191]}
   );
   gpc1_1 gpc1_1_2184(
      {stage064[51]},
      {stage064[192]}
   );
   gpc1_1 gpc1_1_2185(
      {stage064[52]},
      {stage064[193]}
   );
   gpc1_1 gpc1_1_2186(
      {stage064[53]},
      {stage064[194]}
   );
   gpc1_1 gpc1_1_2187(
      {stage064[54]},
      {stage064[195]}
   );
   gpc1_1 gpc1_1_2188(
      {stage064[55]},
      {stage064[196]}
   );
   gpc1_1 gpc1_1_2189(
      {stage064[56]},
      {stage064[197]}
   );
   gpc606_5 gpc606_5_2190(
      {stage064[57], stage064[58], stage064[59], stage064[60], stage064[61], stage064[62]},
      {stage066[0], stage066[1], stage066[2], stage066[3], stage066[4], stage066[5]},
      {stage068[128], stage067[135], stage066[139], stage065[152], stage064[198]}
   );
   gpc606_5 gpc606_5_2191(
      {stage064[63], stage064[64], stage064[65], stage064[66], stage064[67], stage064[68]},
      {stage066[6], stage066[7], stage066[8], stage066[9], stage066[10], stage066[11]},
      {stage068[129], stage067[136], stage066[140], stage065[153], stage064[199]}
   );
   gpc606_5 gpc606_5_2192(
      {stage064[69], stage064[70], stage064[71], stage064[72], stage064[73], stage064[74]},
      {stage066[12], stage066[13], stage066[14], stage066[15], stage066[16], stage066[17]},
      {stage068[130], stage067[137], stage066[141], stage065[154], stage064[200]}
   );
   gpc606_5 gpc606_5_2193(
      {stage064[75], stage064[76], stage064[77], stage064[78], stage064[79], stage064[80]},
      {stage066[18], stage066[19], stage066[20], stage066[21], stage066[22], stage066[23]},
      {stage068[131], stage067[138], stage066[142], stage065[155], stage064[201]}
   );
   gpc606_5 gpc606_5_2194(
      {stage064[81], stage064[82], stage064[83], stage064[84], stage064[85], stage064[86]},
      {stage066[24], stage066[25], stage066[26], stage066[27], stage066[28], stage066[29]},
      {stage068[132], stage067[139], stage066[143], stage065[156], stage064[202]}
   );
   gpc606_5 gpc606_5_2195(
      {stage064[87], stage064[88], stage064[89], stage064[90], stage064[91], stage064[92]},
      {stage066[30], stage066[31], stage066[32], stage066[33], stage066[34], stage066[35]},
      {stage068[133], stage067[140], stage066[144], stage065[157], stage064[203]}
   );
   gpc615_5 gpc615_5_2196(
      {stage064[93], stage064[94], stage064[95], stage064[96], stage064[97]},
      {stage065[42]},
      {stage066[36], stage066[37], stage066[38], stage066[39], stage066[40], stage066[41]},
      {stage068[134], stage067[141], stage066[145], stage065[158], stage064[204]}
   );
   gpc615_5 gpc615_5_2197(
      {stage064[98], stage064[99], stage064[100], stage064[101], stage064[102]},
      {stage065[43]},
      {stage066[42], stage066[43], stage066[44], stage066[45], stage066[46], stage066[47]},
      {stage068[135], stage067[142], stage066[146], stage065[159], stage064[205]}
   );
   gpc615_5 gpc615_5_2198(
      {stage064[103], stage064[104], stage064[105], stage064[106], stage064[107]},
      {stage065[44]},
      {stage066[48], stage066[49], stage066[50], stage066[51], stage066[52], stage066[53]},
      {stage068[136], stage067[143], stage066[147], stage065[160], stage064[206]}
   );
   gpc615_5 gpc615_5_2199(
      {stage064[108], stage064[109], stage064[110], stage064[111], stage064[112]},
      {stage065[45]},
      {stage066[54], stage066[55], stage066[56], stage066[57], stage066[58], stage066[59]},
      {stage068[137], stage067[144], stage066[148], stage065[161], stage064[207]}
   );
   gpc615_5 gpc615_5_2200(
      {stage064[113], stage064[114], stage064[115], stage064[116], stage064[117]},
      {stage065[46]},
      {stage066[60], stage066[61], stage066[62], stage066[63], stage066[64], stage066[65]},
      {stage068[138], stage067[145], stage066[149], stage065[162], stage064[208]}
   );
   gpc615_5 gpc615_5_2201(
      {stage064[118], stage064[119], stage064[120], stage064[121], stage064[122]},
      {stage065[47]},
      {stage066[66], stage066[67], stage066[68], stage066[69], stage066[70], stage066[71]},
      {stage068[139], stage067[146], stage066[150], stage065[163], stage064[209]}
   );
   gpc615_5 gpc615_5_2202(
      {stage064[123], stage064[124], stage064[125], stage064[126], stage064[127]},
      {stage065[48]},
      {stage066[72], stage066[73], stage066[74], stage066[75], stage066[76], stage066[77]},
      {stage068[140], stage067[147], stage066[151], stage065[164], stage064[210]}
   );
   gpc1_1 gpc1_1_2203(
      {stage065[49]},
      {stage065[165]}
   );
   gpc1_1 gpc1_1_2204(
      {stage065[50]},
      {stage065[166]}
   );
   gpc1_1 gpc1_1_2205(
      {stage065[51]},
      {stage065[167]}
   );
   gpc1_1 gpc1_1_2206(
      {stage065[52]},
      {stage065[168]}
   );
   gpc1_1 gpc1_1_2207(
      {stage065[53]},
      {stage065[169]}
   );
   gpc1_1 gpc1_1_2208(
      {stage065[54]},
      {stage065[170]}
   );
   gpc1_1 gpc1_1_2209(
      {stage065[55]},
      {stage065[171]}
   );
   gpc1_1 gpc1_1_2210(
      {stage065[56]},
      {stage065[172]}
   );
   gpc1_1 gpc1_1_2211(
      {stage065[57]},
      {stage065[173]}
   );
   gpc1_1 gpc1_1_2212(
      {stage065[58]},
      {stage065[174]}
   );
   gpc1_1 gpc1_1_2213(
      {stage065[59]},
      {stage065[175]}
   );
   gpc1_1 gpc1_1_2214(
      {stage065[60]},
      {stage065[176]}
   );
   gpc1_1 gpc1_1_2215(
      {stage065[61]},
      {stage065[177]}
   );
   gpc1_1 gpc1_1_2216(
      {stage065[62]},
      {stage065[178]}
   );
   gpc1_1 gpc1_1_2217(
      {stage065[63]},
      {stage065[179]}
   );
   gpc1_1 gpc1_1_2218(
      {stage065[64]},
      {stage065[180]}
   );
   gpc1_1 gpc1_1_2219(
      {stage065[65]},
      {stage065[181]}
   );
   gpc1_1 gpc1_1_2220(
      {stage065[66]},
      {stage065[182]}
   );
   gpc1_1 gpc1_1_2221(
      {stage065[67]},
      {stage065[183]}
   );
   gpc1_1 gpc1_1_2222(
      {stage065[68]},
      {stage065[184]}
   );
   gpc1_1 gpc1_1_2223(
      {stage065[69]},
      {stage065[185]}
   );
   gpc1_1 gpc1_1_2224(
      {stage065[70]},
      {stage065[186]}
   );
   gpc1_1 gpc1_1_2225(
      {stage065[71]},
      {stage065[187]}
   );
   gpc1_1 gpc1_1_2226(
      {stage065[72]},
      {stage065[188]}
   );
   gpc1_1 gpc1_1_2227(
      {stage065[73]},
      {stage065[189]}
   );
   gpc606_5 gpc606_5_2228(
      {stage065[74], stage065[75], stage065[76], stage065[77], stage065[78], stage065[79]},
      {stage067[0], stage067[1], stage067[2], stage067[3], stage067[4], stage067[5]},
      {stage069[128], stage068[141], stage067[148], stage066[152], stage065[190]}
   );
   gpc606_5 gpc606_5_2229(
      {stage065[80], stage065[81], stage065[82], stage065[83], stage065[84], stage065[85]},
      {stage067[6], stage067[7], stage067[8], stage067[9], stage067[10], stage067[11]},
      {stage069[129], stage068[142], stage067[149], stage066[153], stage065[191]}
   );
   gpc606_5 gpc606_5_2230(
      {stage065[86], stage065[87], stage065[88], stage065[89], stage065[90], stage065[91]},
      {stage067[12], stage067[13], stage067[14], stage067[15], stage067[16], stage067[17]},
      {stage069[130], stage068[143], stage067[150], stage066[154], stage065[192]}
   );
   gpc606_5 gpc606_5_2231(
      {stage065[92], stage065[93], stage065[94], stage065[95], stage065[96], stage065[97]},
      {stage067[18], stage067[19], stage067[20], stage067[21], stage067[22], stage067[23]},
      {stage069[131], stage068[144], stage067[151], stage066[155], stage065[193]}
   );
   gpc606_5 gpc606_5_2232(
      {stage065[98], stage065[99], stage065[100], stage065[101], stage065[102], stage065[103]},
      {stage067[24], stage067[25], stage067[26], stage067[27], stage067[28], stage067[29]},
      {stage069[132], stage068[145], stage067[152], stage066[156], stage065[194]}
   );
   gpc606_5 gpc606_5_2233(
      {stage065[104], stage065[105], stage065[106], stage065[107], stage065[108], stage065[109]},
      {stage067[30], stage067[31], stage067[32], stage067[33], stage067[34], stage067[35]},
      {stage069[133], stage068[146], stage067[153], stage066[157], stage065[195]}
   );
   gpc606_5 gpc606_5_2234(
      {stage065[110], stage065[111], stage065[112], stage065[113], stage065[114], stage065[115]},
      {stage067[36], stage067[37], stage067[38], stage067[39], stage067[40], stage067[41]},
      {stage069[134], stage068[147], stage067[154], stage066[158], stage065[196]}
   );
   gpc606_5 gpc606_5_2235(
      {stage065[116], stage065[117], stage065[118], stage065[119], stage065[120], stage065[121]},
      {stage067[42], stage067[43], stage067[44], stage067[45], stage067[46], stage067[47]},
      {stage069[135], stage068[148], stage067[155], stage066[159], stage065[197]}
   );
   gpc606_5 gpc606_5_2236(
      {stage065[122], stage065[123], stage065[124], stage065[125], stage065[126], stage065[127]},
      {stage067[48], stage067[49], stage067[50], stage067[51], stage067[52], stage067[53]},
      {stage069[136], stage068[149], stage067[156], stage066[160], stage065[198]}
   );
   gpc1_1 gpc1_1_2237(
      {stage066[78]},
      {stage066[161]}
   );
   gpc1_1 gpc1_1_2238(
      {stage066[79]},
      {stage066[162]}
   );
   gpc1_1 gpc1_1_2239(
      {stage066[80]},
      {stage066[163]}
   );
   gpc1_1 gpc1_1_2240(
      {stage066[81]},
      {stage066[164]}
   );
   gpc1_1 gpc1_1_2241(
      {stage066[82]},
      {stage066[165]}
   );
   gpc1_1 gpc1_1_2242(
      {stage066[83]},
      {stage066[166]}
   );
   gpc1_1 gpc1_1_2243(
      {stage066[84]},
      {stage066[167]}
   );
   gpc1_1 gpc1_1_2244(
      {stage066[85]},
      {stage066[168]}
   );
   gpc1_1 gpc1_1_2245(
      {stage066[86]},
      {stage066[169]}
   );
   gpc1_1 gpc1_1_2246(
      {stage066[87]},
      {stage066[170]}
   );
   gpc1_1 gpc1_1_2247(
      {stage066[88]},
      {stage066[171]}
   );
   gpc1_1 gpc1_1_2248(
      {stage066[89]},
      {stage066[172]}
   );
   gpc1_1 gpc1_1_2249(
      {stage066[90]},
      {stage066[173]}
   );
   gpc1_1 gpc1_1_2250(
      {stage066[91]},
      {stage066[174]}
   );
   gpc1_1 gpc1_1_2251(
      {stage066[92]},
      {stage066[175]}
   );
   gpc1_1 gpc1_1_2252(
      {stage066[93]},
      {stage066[176]}
   );
   gpc1_1 gpc1_1_2253(
      {stage066[94]},
      {stage066[177]}
   );
   gpc1_1 gpc1_1_2254(
      {stage066[95]},
      {stage066[178]}
   );
   gpc1_1 gpc1_1_2255(
      {stage066[96]},
      {stage066[179]}
   );
   gpc1_1 gpc1_1_2256(
      {stage066[97]},
      {stage066[180]}
   );
   gpc1_1 gpc1_1_2257(
      {stage066[98]},
      {stage066[181]}
   );
   gpc1_1 gpc1_1_2258(
      {stage066[99]},
      {stage066[182]}
   );
   gpc1_1 gpc1_1_2259(
      {stage066[100]},
      {stage066[183]}
   );
   gpc1_1 gpc1_1_2260(
      {stage066[101]},
      {stage066[184]}
   );
   gpc1_1 gpc1_1_2261(
      {stage066[102]},
      {stage066[185]}
   );
   gpc1_1 gpc1_1_2262(
      {stage066[103]},
      {stage066[186]}
   );
   gpc1_1 gpc1_1_2263(
      {stage066[104]},
      {stage066[187]}
   );
   gpc1_1 gpc1_1_2264(
      {stage066[105]},
      {stage066[188]}
   );
   gpc1_1 gpc1_1_2265(
      {stage066[106]},
      {stage066[189]}
   );
   gpc1_1 gpc1_1_2266(
      {stage066[107]},
      {stage066[190]}
   );
   gpc1_1 gpc1_1_2267(
      {stage066[108]},
      {stage066[191]}
   );
   gpc1_1 gpc1_1_2268(
      {stage066[109]},
      {stage066[192]}
   );
   gpc1_1 gpc1_1_2269(
      {stage066[110]},
      {stage066[193]}
   );
   gpc1_1 gpc1_1_2270(
      {stage066[111]},
      {stage066[194]}
   );
   gpc1_1 gpc1_1_2271(
      {stage066[112]},
      {stage066[195]}
   );
   gpc1_1 gpc1_1_2272(
      {stage066[113]},
      {stage066[196]}
   );
   gpc1_1 gpc1_1_2273(
      {stage066[114]},
      {stage066[197]}
   );
   gpc1_1 gpc1_1_2274(
      {stage066[115]},
      {stage066[198]}
   );
   gpc1_1 gpc1_1_2275(
      {stage066[116]},
      {stage066[199]}
   );
   gpc1_1 gpc1_1_2276(
      {stage066[117]},
      {stage066[200]}
   );
   gpc1_1 gpc1_1_2277(
      {stage066[118]},
      {stage066[201]}
   );
   gpc1_1 gpc1_1_2278(
      {stage066[119]},
      {stage066[202]}
   );
   gpc1_1 gpc1_1_2279(
      {stage066[120]},
      {stage066[203]}
   );
   gpc1_1 gpc1_1_2280(
      {stage066[121]},
      {stage066[204]}
   );
   gpc1_1 gpc1_1_2281(
      {stage066[122]},
      {stage066[205]}
   );
   gpc1_1 gpc1_1_2282(
      {stage066[123]},
      {stage066[206]}
   );
   gpc1_1 gpc1_1_2283(
      {stage066[124]},
      {stage066[207]}
   );
   gpc1_1 gpc1_1_2284(
      {stage066[125]},
      {stage066[208]}
   );
   gpc1_1 gpc1_1_2285(
      {stage066[126]},
      {stage066[209]}
   );
   gpc1_1 gpc1_1_2286(
      {stage066[127]},
      {stage066[210]}
   );
   gpc1_1 gpc1_1_2287(
      {stage067[54]},
      {stage067[157]}
   );
   gpc1_1 gpc1_1_2288(
      {stage067[55]},
      {stage067[158]}
   );
   gpc1_1 gpc1_1_2289(
      {stage067[56]},
      {stage067[159]}
   );
   gpc1_1 gpc1_1_2290(
      {stage067[57]},
      {stage067[160]}
   );
   gpc1_1 gpc1_1_2291(
      {stage067[58]},
      {stage067[161]}
   );
   gpc1_1 gpc1_1_2292(
      {stage067[59]},
      {stage067[162]}
   );
   gpc1_1 gpc1_1_2293(
      {stage067[60]},
      {stage067[163]}
   );
   gpc1_1 gpc1_1_2294(
      {stage067[61]},
      {stage067[164]}
   );
   gpc1_1 gpc1_1_2295(
      {stage067[62]},
      {stage067[165]}
   );
   gpc1_1 gpc1_1_2296(
      {stage067[63]},
      {stage067[166]}
   );
   gpc1_1 gpc1_1_2297(
      {stage067[64]},
      {stage067[167]}
   );
   gpc1_1 gpc1_1_2298(
      {stage067[65]},
      {stage067[168]}
   );
   gpc1_1 gpc1_1_2299(
      {stage067[66]},
      {stage067[169]}
   );
   gpc1_1 gpc1_1_2300(
      {stage067[67]},
      {stage067[170]}
   );
   gpc1_1 gpc1_1_2301(
      {stage067[68]},
      {stage067[171]}
   );
   gpc1_1 gpc1_1_2302(
      {stage067[69]},
      {stage067[172]}
   );
   gpc1_1 gpc1_1_2303(
      {stage067[70]},
      {stage067[173]}
   );
   gpc1_1 gpc1_1_2304(
      {stage067[71]},
      {stage067[174]}
   );
   gpc1_1 gpc1_1_2305(
      {stage067[72]},
      {stage067[175]}
   );
   gpc1_1 gpc1_1_2306(
      {stage067[73]},
      {stage067[176]}
   );
   gpc1_1 gpc1_1_2307(
      {stage067[74]},
      {stage067[177]}
   );
   gpc1_1 gpc1_1_2308(
      {stage067[75]},
      {stage067[178]}
   );
   gpc1_1 gpc1_1_2309(
      {stage067[76]},
      {stage067[179]}
   );
   gpc1_1 gpc1_1_2310(
      {stage067[77]},
      {stage067[180]}
   );
   gpc1_1 gpc1_1_2311(
      {stage067[78]},
      {stage067[181]}
   );
   gpc1_1 gpc1_1_2312(
      {stage067[79]},
      {stage067[182]}
   );
   gpc1_1 gpc1_1_2313(
      {stage067[80]},
      {stage067[183]}
   );
   gpc1_1 gpc1_1_2314(
      {stage067[81]},
      {stage067[184]}
   );
   gpc1_1 gpc1_1_2315(
      {stage067[82]},
      {stage067[185]}
   );
   gpc1_1 gpc1_1_2316(
      {stage067[83]},
      {stage067[186]}
   );
   gpc1_1 gpc1_1_2317(
      {stage067[84]},
      {stage067[187]}
   );
   gpc1_1 gpc1_1_2318(
      {stage067[85]},
      {stage067[188]}
   );
   gpc1_1 gpc1_1_2319(
      {stage067[86]},
      {stage067[189]}
   );
   gpc1_1 gpc1_1_2320(
      {stage067[87]},
      {stage067[190]}
   );
   gpc1_1 gpc1_1_2321(
      {stage067[88]},
      {stage067[191]}
   );
   gpc1_1 gpc1_1_2322(
      {stage067[89]},
      {stage067[192]}
   );
   gpc1_1 gpc1_1_2323(
      {stage067[90]},
      {stage067[193]}
   );
   gpc1_1 gpc1_1_2324(
      {stage067[91]},
      {stage067[194]}
   );
   gpc1_1 gpc1_1_2325(
      {stage067[92]},
      {stage067[195]}
   );
   gpc1_1 gpc1_1_2326(
      {stage067[93]},
      {stage067[196]}
   );
   gpc1_1 gpc1_1_2327(
      {stage067[94]},
      {stage067[197]}
   );
   gpc1_1 gpc1_1_2328(
      {stage067[95]},
      {stage067[198]}
   );
   gpc1_1 gpc1_1_2329(
      {stage067[96]},
      {stage067[199]}
   );
   gpc1_1 gpc1_1_2330(
      {stage067[97]},
      {stage067[200]}
   );
   gpc1_1 gpc1_1_2331(
      {stage067[98]},
      {stage067[201]}
   );
   gpc1_1 gpc1_1_2332(
      {stage067[99]},
      {stage067[202]}
   );
   gpc1_1 gpc1_1_2333(
      {stage067[100]},
      {stage067[203]}
   );
   gpc1_1 gpc1_1_2334(
      {stage067[101]},
      {stage067[204]}
   );
   gpc1_1 gpc1_1_2335(
      {stage067[102]},
      {stage067[205]}
   );
   gpc1_1 gpc1_1_2336(
      {stage067[103]},
      {stage067[206]}
   );
   gpc1_1 gpc1_1_2337(
      {stage067[104]},
      {stage067[207]}
   );
   gpc1_1 gpc1_1_2338(
      {stage067[105]},
      {stage067[208]}
   );
   gpc606_5 gpc606_5_2339(
      {stage067[106], stage067[107], stage067[108], stage067[109], stage067[110], stage067[111]},
      {stage069[0], stage069[1], stage069[2], stage069[3], stage069[4], stage069[5]},
      {stage071[128], stage070[128], stage069[137], stage068[150], stage067[209]}
   );
   gpc606_5 gpc606_5_2340(
      {stage067[112], stage067[113], stage067[114], stage067[115], stage067[116], stage067[117]},
      {stage069[6], stage069[7], stage069[8], stage069[9], stage069[10], stage069[11]},
      {stage071[129], stage070[129], stage069[138], stage068[151], stage067[210]}
   );
   gpc615_5 gpc615_5_2341(
      {stage067[118], stage067[119], stage067[120], stage067[121], stage067[122]},
      {stage068[0]},
      {stage069[12], stage069[13], stage069[14], stage069[15], stage069[16], stage069[17]},
      {stage071[130], stage070[130], stage069[139], stage068[152], stage067[211]}
   );
   gpc1325_5 gpc1325_5_2342(
      {stage067[123], stage067[124], stage067[125], stage067[126], stage067[127]},
      {stage068[1], stage068[2]},
      {stage069[18], stage069[19], stage069[20]},
      {stage070[0]},
      {stage071[131], stage070[131], stage069[140], stage068[153], stage067[212]}
   );
   gpc1_1 gpc1_1_2343(
      {stage068[3]},
      {stage068[154]}
   );
   gpc1_1 gpc1_1_2344(
      {stage068[4]},
      {stage068[155]}
   );
   gpc1_1 gpc1_1_2345(
      {stage068[5]},
      {stage068[156]}
   );
   gpc1_1 gpc1_1_2346(
      {stage068[6]},
      {stage068[157]}
   );
   gpc1_1 gpc1_1_2347(
      {stage068[7]},
      {stage068[158]}
   );
   gpc1_1 gpc1_1_2348(
      {stage068[8]},
      {stage068[159]}
   );
   gpc1_1 gpc1_1_2349(
      {stage068[9]},
      {stage068[160]}
   );
   gpc1_1 gpc1_1_2350(
      {stage068[10]},
      {stage068[161]}
   );
   gpc1_1 gpc1_1_2351(
      {stage068[11]},
      {stage068[162]}
   );
   gpc1_1 gpc1_1_2352(
      {stage068[12]},
      {stage068[163]}
   );
   gpc1_1 gpc1_1_2353(
      {stage068[13]},
      {stage068[164]}
   );
   gpc1_1 gpc1_1_2354(
      {stage068[14]},
      {stage068[165]}
   );
   gpc1_1 gpc1_1_2355(
      {stage068[15]},
      {stage068[166]}
   );
   gpc1_1 gpc1_1_2356(
      {stage068[16]},
      {stage068[167]}
   );
   gpc1_1 gpc1_1_2357(
      {stage068[17]},
      {stage068[168]}
   );
   gpc1_1 gpc1_1_2358(
      {stage068[18]},
      {stage068[169]}
   );
   gpc1_1 gpc1_1_2359(
      {stage068[19]},
      {stage068[170]}
   );
   gpc1_1 gpc1_1_2360(
      {stage068[20]},
      {stage068[171]}
   );
   gpc1_1 gpc1_1_2361(
      {stage068[21]},
      {stage068[172]}
   );
   gpc1_1 gpc1_1_2362(
      {stage068[22]},
      {stage068[173]}
   );
   gpc1_1 gpc1_1_2363(
      {stage068[23]},
      {stage068[174]}
   );
   gpc1_1 gpc1_1_2364(
      {stage068[24]},
      {stage068[175]}
   );
   gpc1_1 gpc1_1_2365(
      {stage068[25]},
      {stage068[176]}
   );
   gpc1_1 gpc1_1_2366(
      {stage068[26]},
      {stage068[177]}
   );
   gpc1_1 gpc1_1_2367(
      {stage068[27]},
      {stage068[178]}
   );
   gpc1_1 gpc1_1_2368(
      {stage068[28]},
      {stage068[179]}
   );
   gpc1_1 gpc1_1_2369(
      {stage068[29]},
      {stage068[180]}
   );
   gpc1_1 gpc1_1_2370(
      {stage068[30]},
      {stage068[181]}
   );
   gpc1_1 gpc1_1_2371(
      {stage068[31]},
      {stage068[182]}
   );
   gpc1_1 gpc1_1_2372(
      {stage068[32]},
      {stage068[183]}
   );
   gpc1_1 gpc1_1_2373(
      {stage068[33]},
      {stage068[184]}
   );
   gpc1_1 gpc1_1_2374(
      {stage068[34]},
      {stage068[185]}
   );
   gpc1_1 gpc1_1_2375(
      {stage068[35]},
      {stage068[186]}
   );
   gpc1_1 gpc1_1_2376(
      {stage068[36]},
      {stage068[187]}
   );
   gpc1_1 gpc1_1_2377(
      {stage068[37]},
      {stage068[188]}
   );
   gpc1_1 gpc1_1_2378(
      {stage068[38]},
      {stage068[189]}
   );
   gpc1_1 gpc1_1_2379(
      {stage068[39]},
      {stage068[190]}
   );
   gpc1_1 gpc1_1_2380(
      {stage068[40]},
      {stage068[191]}
   );
   gpc1_1 gpc1_1_2381(
      {stage068[41]},
      {stage068[192]}
   );
   gpc1_1 gpc1_1_2382(
      {stage068[42]},
      {stage068[193]}
   );
   gpc1_1 gpc1_1_2383(
      {stage068[43]},
      {stage068[194]}
   );
   gpc1_1 gpc1_1_2384(
      {stage068[44]},
      {stage068[195]}
   );
   gpc606_5 gpc606_5_2385(
      {stage068[45], stage068[46], stage068[47], stage068[48], stage068[49], stage068[50]},
      {stage070[1], stage070[2], stage070[3], stage070[4], stage070[5], stage070[6]},
      {stage072[128], stage071[132], stage070[132], stage069[141], stage068[196]}
   );
   gpc606_5 gpc606_5_2386(
      {stage068[51], stage068[52], stage068[53], stage068[54], stage068[55], stage068[56]},
      {stage070[7], stage070[8], stage070[9], stage070[10], stage070[11], stage070[12]},
      {stage072[129], stage071[133], stage070[133], stage069[142], stage068[197]}
   );
   gpc606_5 gpc606_5_2387(
      {stage068[57], stage068[58], stage068[59], stage068[60], stage068[61], stage068[62]},
      {stage070[13], stage070[14], stage070[15], stage070[16], stage070[17], stage070[18]},
      {stage072[130], stage071[134], stage070[134], stage069[143], stage068[198]}
   );
   gpc606_5 gpc606_5_2388(
      {stage068[63], stage068[64], stage068[65], stage068[66], stage068[67], stage068[68]},
      {stage070[19], stage070[20], stage070[21], stage070[22], stage070[23], stage070[24]},
      {stage072[131], stage071[135], stage070[135], stage069[144], stage068[199]}
   );
   gpc606_5 gpc606_5_2389(
      {stage068[69], stage068[70], stage068[71], stage068[72], stage068[73], stage068[74]},
      {stage070[25], stage070[26], stage070[27], stage070[28], stage070[29], stage070[30]},
      {stage072[132], stage071[136], stage070[136], stage069[145], stage068[200]}
   );
   gpc606_5 gpc606_5_2390(
      {stage068[75], stage068[76], stage068[77], stage068[78], stage068[79], stage068[80]},
      {stage070[31], stage070[32], stage070[33], stage070[34], stage070[35], stage070[36]},
      {stage072[133], stage071[137], stage070[137], stage069[146], stage068[201]}
   );
   gpc606_5 gpc606_5_2391(
      {stage068[81], stage068[82], stage068[83], stage068[84], stage068[85], stage068[86]},
      {stage070[37], stage070[38], stage070[39], stage070[40], stage070[41], stage070[42]},
      {stage072[134], stage071[138], stage070[138], stage069[147], stage068[202]}
   );
   gpc606_5 gpc606_5_2392(
      {stage068[87], stage068[88], stage068[89], stage068[90], stage068[91], stage068[92]},
      {stage070[43], stage070[44], stage070[45], stage070[46], stage070[47], stage070[48]},
      {stage072[135], stage071[139], stage070[139], stage069[148], stage068[203]}
   );
   gpc606_5 gpc606_5_2393(
      {stage068[93], stage068[94], stage068[95], stage068[96], stage068[97], stage068[98]},
      {stage070[49], stage070[50], stage070[51], stage070[52], stage070[53], stage070[54]},
      {stage072[136], stage071[140], stage070[140], stage069[149], stage068[204]}
   );
   gpc606_5 gpc606_5_2394(
      {stage068[99], stage068[100], stage068[101], stage068[102], stage068[103], stage068[104]},
      {stage070[55], stage070[56], stage070[57], stage070[58], stage070[59], stage070[60]},
      {stage072[137], stage071[141], stage070[141], stage069[150], stage068[205]}
   );
   gpc606_5 gpc606_5_2395(
      {stage068[105], stage068[106], stage068[107], stage068[108], stage068[109], stage068[110]},
      {stage070[61], stage070[62], stage070[63], stage070[64], stage070[65], stage070[66]},
      {stage072[138], stage071[142], stage070[142], stage069[151], stage068[206]}
   );
   gpc606_5 gpc606_5_2396(
      {stage068[111], stage068[112], stage068[113], stage068[114], stage068[115], stage068[116]},
      {stage070[67], stage070[68], stage070[69], stage070[70], stage070[71], stage070[72]},
      {stage072[139], stage071[143], stage070[143], stage069[152], stage068[207]}
   );
   gpc606_5 gpc606_5_2397(
      {stage068[117], stage068[118], stage068[119], stage068[120], stage068[121], stage068[122]},
      {stage070[73], stage070[74], stage070[75], stage070[76], stage070[77], stage070[78]},
      {stage072[140], stage071[144], stage070[144], stage069[153], stage068[208]}
   );
   gpc2135_5 gpc2135_5_2398(
      {stage068[123], stage068[124], stage068[125], stage068[126], stage068[127]},
      {stage069[21], stage069[22], stage069[23]},
      {stage070[79]},
      {stage071[0], stage071[1]},
      {stage072[141], stage071[145], stage070[145], stage069[154], stage068[209]}
   );
   gpc1_1 gpc1_1_2399(
      {stage069[24]},
      {stage069[155]}
   );
   gpc1_1 gpc1_1_2400(
      {stage069[25]},
      {stage069[156]}
   );
   gpc1_1 gpc1_1_2401(
      {stage069[26]},
      {stage069[157]}
   );
   gpc1_1 gpc1_1_2402(
      {stage069[27]},
      {stage069[158]}
   );
   gpc1_1 gpc1_1_2403(
      {stage069[28]},
      {stage069[159]}
   );
   gpc1_1 gpc1_1_2404(
      {stage069[29]},
      {stage069[160]}
   );
   gpc1_1 gpc1_1_2405(
      {stage069[30]},
      {stage069[161]}
   );
   gpc1_1 gpc1_1_2406(
      {stage069[31]},
      {stage069[162]}
   );
   gpc1_1 gpc1_1_2407(
      {stage069[32]},
      {stage069[163]}
   );
   gpc1_1 gpc1_1_2408(
      {stage069[33]},
      {stage069[164]}
   );
   gpc1_1 gpc1_1_2409(
      {stage069[34]},
      {stage069[165]}
   );
   gpc1_1 gpc1_1_2410(
      {stage069[35]},
      {stage069[166]}
   );
   gpc1_1 gpc1_1_2411(
      {stage069[36]},
      {stage069[167]}
   );
   gpc7_3 gpc7_3_2412(
      {stage069[37], stage069[38], stage069[39], stage069[40], stage069[41], stage069[42], stage069[43]},
      {stage071[146], stage070[146], stage069[168]}
   );
   gpc606_5 gpc606_5_2413(
      {stage069[44], stage069[45], stage069[46], stage069[47], stage069[48], stage069[49]},
      {stage071[2], stage071[3], stage071[4], stage071[5], stage071[6], stage071[7]},
      {stage073[128], stage072[142], stage071[147], stage070[147], stage069[169]}
   );
   gpc606_5 gpc606_5_2414(
      {stage069[50], stage069[51], stage069[52], stage069[53], stage069[54], stage069[55]},
      {stage071[8], stage071[9], stage071[10], stage071[11], stage071[12], stage071[13]},
      {stage073[129], stage072[143], stage071[148], stage070[148], stage069[170]}
   );
   gpc606_5 gpc606_5_2415(
      {stage069[56], stage069[57], stage069[58], stage069[59], stage069[60], stage069[61]},
      {stage071[14], stage071[15], stage071[16], stage071[17], stage071[18], stage071[19]},
      {stage073[130], stage072[144], stage071[149], stage070[149], stage069[171]}
   );
   gpc606_5 gpc606_5_2416(
      {stage069[62], stage069[63], stage069[64], stage069[65], stage069[66], stage069[67]},
      {stage071[20], stage071[21], stage071[22], stage071[23], stage071[24], stage071[25]},
      {stage073[131], stage072[145], stage071[150], stage070[150], stage069[172]}
   );
   gpc606_5 gpc606_5_2417(
      {stage069[68], stage069[69], stage069[70], stage069[71], stage069[72], stage069[73]},
      {stage071[26], stage071[27], stage071[28], stage071[29], stage071[30], stage071[31]},
      {stage073[132], stage072[146], stage071[151], stage070[151], stage069[173]}
   );
   gpc606_5 gpc606_5_2418(
      {stage069[74], stage069[75], stage069[76], stage069[77], stage069[78], stage069[79]},
      {stage071[32], stage071[33], stage071[34], stage071[35], stage071[36], stage071[37]},
      {stage073[133], stage072[147], stage071[152], stage070[152], stage069[174]}
   );
   gpc606_5 gpc606_5_2419(
      {stage069[80], stage069[81], stage069[82], stage069[83], stage069[84], stage069[85]},
      {stage071[38], stage071[39], stage071[40], stage071[41], stage071[42], stage071[43]},
      {stage073[134], stage072[148], stage071[153], stage070[153], stage069[175]}
   );
   gpc606_5 gpc606_5_2420(
      {stage069[86], stage069[87], stage069[88], stage069[89], stage069[90], stage069[91]},
      {stage071[44], stage071[45], stage071[46], stage071[47], stage071[48], stage071[49]},
      {stage073[135], stage072[149], stage071[154], stage070[154], stage069[176]}
   );
   gpc606_5 gpc606_5_2421(
      {stage069[92], stage069[93], stage069[94], stage069[95], stage069[96], stage069[97]},
      {stage071[50], stage071[51], stage071[52], stage071[53], stage071[54], stage071[55]},
      {stage073[136], stage072[150], stage071[155], stage070[155], stage069[177]}
   );
   gpc606_5 gpc606_5_2422(
      {stage069[98], stage069[99], stage069[100], stage069[101], stage069[102], stage069[103]},
      {stage071[56], stage071[57], stage071[58], stage071[59], stage071[60], stage071[61]},
      {stage073[137], stage072[151], stage071[156], stage070[156], stage069[178]}
   );
   gpc606_5 gpc606_5_2423(
      {stage069[104], stage069[105], stage069[106], stage069[107], stage069[108], stage069[109]},
      {stage071[62], stage071[63], stage071[64], stage071[65], stage071[66], stage071[67]},
      {stage073[138], stage072[152], stage071[157], stage070[157], stage069[179]}
   );
   gpc606_5 gpc606_5_2424(
      {stage069[110], stage069[111], stage069[112], stage069[113], stage069[114], stage069[115]},
      {stage071[68], stage071[69], stage071[70], stage071[71], stage071[72], stage071[73]},
      {stage073[139], stage072[153], stage071[158], stage070[158], stage069[180]}
   );
   gpc606_5 gpc606_5_2425(
      {stage069[116], stage069[117], stage069[118], stage069[119], stage069[120], stage069[121]},
      {stage071[74], stage071[75], stage071[76], stage071[77], stage071[78], stage071[79]},
      {stage073[140], stage072[154], stage071[159], stage070[159], stage069[181]}
   );
   gpc606_5 gpc606_5_2426(
      {stage069[122], stage069[123], stage069[124], stage069[125], stage069[126], stage069[127]},
      {stage071[80], stage071[81], stage071[82], stage071[83], stage071[84], stage071[85]},
      {stage073[141], stage072[155], stage071[160], stage070[160], stage069[182]}
   );
   gpc1_1 gpc1_1_2427(
      {stage070[80]},
      {stage070[161]}
   );
   gpc1_1 gpc1_1_2428(
      {stage070[81]},
      {stage070[162]}
   );
   gpc1_1 gpc1_1_2429(
      {stage070[82]},
      {stage070[163]}
   );
   gpc1_1 gpc1_1_2430(
      {stage070[83]},
      {stage070[164]}
   );
   gpc1_1 gpc1_1_2431(
      {stage070[84]},
      {stage070[165]}
   );
   gpc1_1 gpc1_1_2432(
      {stage070[85]},
      {stage070[166]}
   );
   gpc1_1 gpc1_1_2433(
      {stage070[86]},
      {stage070[167]}
   );
   gpc1_1 gpc1_1_2434(
      {stage070[87]},
      {stage070[168]}
   );
   gpc1_1 gpc1_1_2435(
      {stage070[88]},
      {stage070[169]}
   );
   gpc1_1 gpc1_1_2436(
      {stage070[89]},
      {stage070[170]}
   );
   gpc1_1 gpc1_1_2437(
      {stage070[90]},
      {stage070[171]}
   );
   gpc1_1 gpc1_1_2438(
      {stage070[91]},
      {stage070[172]}
   );
   gpc1_1 gpc1_1_2439(
      {stage070[92]},
      {stage070[173]}
   );
   gpc1_1 gpc1_1_2440(
      {stage070[93]},
      {stage070[174]}
   );
   gpc1_1 gpc1_1_2441(
      {stage070[94]},
      {stage070[175]}
   );
   gpc1_1 gpc1_1_2442(
      {stage070[95]},
      {stage070[176]}
   );
   gpc1_1 gpc1_1_2443(
      {stage070[96]},
      {stage070[177]}
   );
   gpc1_1 gpc1_1_2444(
      {stage070[97]},
      {stage070[178]}
   );
   gpc1_1 gpc1_1_2445(
      {stage070[98]},
      {stage070[179]}
   );
   gpc1_1 gpc1_1_2446(
      {stage070[99]},
      {stage070[180]}
   );
   gpc1_1 gpc1_1_2447(
      {stage070[100]},
      {stage070[181]}
   );
   gpc1_1 gpc1_1_2448(
      {stage070[101]},
      {stage070[182]}
   );
   gpc1_1 gpc1_1_2449(
      {stage070[102]},
      {stage070[183]}
   );
   gpc615_5 gpc615_5_2450(
      {stage070[103], stage070[104], stage070[105], stage070[106], stage070[107]},
      {stage071[86]},
      {stage072[0], stage072[1], stage072[2], stage072[3], stage072[4], stage072[5]},
      {stage074[128], stage073[142], stage072[156], stage071[161], stage070[184]}
   );
   gpc615_5 gpc615_5_2451(
      {stage070[108], stage070[109], stage070[110], stage070[111], stage070[112]},
      {stage071[87]},
      {stage072[6], stage072[7], stage072[8], stage072[9], stage072[10], stage072[11]},
      {stage074[129], stage073[143], stage072[157], stage071[162], stage070[185]}
   );
   gpc615_5 gpc615_5_2452(
      {stage070[113], stage070[114], stage070[115], stage070[116], stage070[117]},
      {stage071[88]},
      {stage072[12], stage072[13], stage072[14], stage072[15], stage072[16], stage072[17]},
      {stage074[130], stage073[144], stage072[158], stage071[163], stage070[186]}
   );
   gpc615_5 gpc615_5_2453(
      {stage070[118], stage070[119], stage070[120], stage070[121], stage070[122]},
      {stage071[89]},
      {stage072[18], stage072[19], stage072[20], stage072[21], stage072[22], stage072[23]},
      {stage074[131], stage073[145], stage072[159], stage071[164], stage070[187]}
   );
   gpc615_5 gpc615_5_2454(
      {stage070[123], stage070[124], stage070[125], stage070[126], stage070[127]},
      {stage071[90]},
      {stage072[24], stage072[25], stage072[26], stage072[27], stage072[28], stage072[29]},
      {stage074[132], stage073[146], stage072[160], stage071[165], stage070[188]}
   );
   gpc1_1 gpc1_1_2455(
      {stage071[91]},
      {stage071[166]}
   );
   gpc1_1 gpc1_1_2456(
      {stage071[92]},
      {stage071[167]}
   );
   gpc1_1 gpc1_1_2457(
      {stage071[93]},
      {stage071[168]}
   );
   gpc1_1 gpc1_1_2458(
      {stage071[94]},
      {stage071[169]}
   );
   gpc1_1 gpc1_1_2459(
      {stage071[95]},
      {stage071[170]}
   );
   gpc1_1 gpc1_1_2460(
      {stage071[96]},
      {stage071[171]}
   );
   gpc1_1 gpc1_1_2461(
      {stage071[97]},
      {stage071[172]}
   );
   gpc1_1 gpc1_1_2462(
      {stage071[98]},
      {stage071[173]}
   );
   gpc1_1 gpc1_1_2463(
      {stage071[99]},
      {stage071[174]}
   );
   gpc1_1 gpc1_1_2464(
      {stage071[100]},
      {stage071[175]}
   );
   gpc1_1 gpc1_1_2465(
      {stage071[101]},
      {stage071[176]}
   );
   gpc1_1 gpc1_1_2466(
      {stage071[102]},
      {stage071[177]}
   );
   gpc1_1 gpc1_1_2467(
      {stage071[103]},
      {stage071[178]}
   );
   gpc1_1 gpc1_1_2468(
      {stage071[104]},
      {stage071[179]}
   );
   gpc1_1 gpc1_1_2469(
      {stage071[105]},
      {stage071[180]}
   );
   gpc1_1 gpc1_1_2470(
      {stage071[106]},
      {stage071[181]}
   );
   gpc1_1 gpc1_1_2471(
      {stage071[107]},
      {stage071[182]}
   );
   gpc1_1 gpc1_1_2472(
      {stage071[108]},
      {stage071[183]}
   );
   gpc1_1 gpc1_1_2473(
      {stage071[109]},
      {stage071[184]}
   );
   gpc606_5 gpc606_5_2474(
      {stage071[110], stage071[111], stage071[112], stage071[113], stage071[114], stage071[115]},
      {stage073[0], stage073[1], stage073[2], stage073[3], stage073[4], stage073[5]},
      {stage075[128], stage074[133], stage073[147], stage072[161], stage071[185]}
   );
   gpc606_5 gpc606_5_2475(
      {stage071[116], stage071[117], stage071[118], stage071[119], stage071[120], stage071[121]},
      {stage073[6], stage073[7], stage073[8], stage073[9], stage073[10], stage073[11]},
      {stage075[129], stage074[134], stage073[148], stage072[162], stage071[186]}
   );
   gpc606_5 gpc606_5_2476(
      {stage071[122], stage071[123], stage071[124], stage071[125], stage071[126], stage071[127]},
      {stage073[12], stage073[13], stage073[14], stage073[15], stage073[16], stage073[17]},
      {stage075[130], stage074[135], stage073[149], stage072[163], stage071[187]}
   );
   gpc1_1 gpc1_1_2477(
      {stage072[30]},
      {stage072[164]}
   );
   gpc1_1 gpc1_1_2478(
      {stage072[31]},
      {stage072[165]}
   );
   gpc1_1 gpc1_1_2479(
      {stage072[32]},
      {stage072[166]}
   );
   gpc1_1 gpc1_1_2480(
      {stage072[33]},
      {stage072[167]}
   );
   gpc1_1 gpc1_1_2481(
      {stage072[34]},
      {stage072[168]}
   );
   gpc1_1 gpc1_1_2482(
      {stage072[35]},
      {stage072[169]}
   );
   gpc1_1 gpc1_1_2483(
      {stage072[36]},
      {stage072[170]}
   );
   gpc1_1 gpc1_1_2484(
      {stage072[37]},
      {stage072[171]}
   );
   gpc1_1 gpc1_1_2485(
      {stage072[38]},
      {stage072[172]}
   );
   gpc1_1 gpc1_1_2486(
      {stage072[39]},
      {stage072[173]}
   );
   gpc1_1 gpc1_1_2487(
      {stage072[40]},
      {stage072[174]}
   );
   gpc1_1 gpc1_1_2488(
      {stage072[41]},
      {stage072[175]}
   );
   gpc1_1 gpc1_1_2489(
      {stage072[42]},
      {stage072[176]}
   );
   gpc1_1 gpc1_1_2490(
      {stage072[43]},
      {stage072[177]}
   );
   gpc1_1 gpc1_1_2491(
      {stage072[44]},
      {stage072[178]}
   );
   gpc1_1 gpc1_1_2492(
      {stage072[45]},
      {stage072[179]}
   );
   gpc1_1 gpc1_1_2493(
      {stage072[46]},
      {stage072[180]}
   );
   gpc1_1 gpc1_1_2494(
      {stage072[47]},
      {stage072[181]}
   );
   gpc1_1 gpc1_1_2495(
      {stage072[48]},
      {stage072[182]}
   );
   gpc1_1 gpc1_1_2496(
      {stage072[49]},
      {stage072[183]}
   );
   gpc1_1 gpc1_1_2497(
      {stage072[50]},
      {stage072[184]}
   );
   gpc1_1 gpc1_1_2498(
      {stage072[51]},
      {stage072[185]}
   );
   gpc1_1 gpc1_1_2499(
      {stage072[52]},
      {stage072[186]}
   );
   gpc1_1 gpc1_1_2500(
      {stage072[53]},
      {stage072[187]}
   );
   gpc1_1 gpc1_1_2501(
      {stage072[54]},
      {stage072[188]}
   );
   gpc1_1 gpc1_1_2502(
      {stage072[55]},
      {stage072[189]}
   );
   gpc1_1 gpc1_1_2503(
      {stage072[56]},
      {stage072[190]}
   );
   gpc1_1 gpc1_1_2504(
      {stage072[57]},
      {stage072[191]}
   );
   gpc1_1 gpc1_1_2505(
      {stage072[58]},
      {stage072[192]}
   );
   gpc1_1 gpc1_1_2506(
      {stage072[59]},
      {stage072[193]}
   );
   gpc1_1 gpc1_1_2507(
      {stage072[60]},
      {stage072[194]}
   );
   gpc1_1 gpc1_1_2508(
      {stage072[61]},
      {stage072[195]}
   );
   gpc1_1 gpc1_1_2509(
      {stage072[62]},
      {stage072[196]}
   );
   gpc1_1 gpc1_1_2510(
      {stage072[63]},
      {stage072[197]}
   );
   gpc1_1 gpc1_1_2511(
      {stage072[64]},
      {stage072[198]}
   );
   gpc1_1 gpc1_1_2512(
      {stage072[65]},
      {stage072[199]}
   );
   gpc1_1 gpc1_1_2513(
      {stage072[66]},
      {stage072[200]}
   );
   gpc1_1 gpc1_1_2514(
      {stage072[67]},
      {stage072[201]}
   );
   gpc1_1 gpc1_1_2515(
      {stage072[68]},
      {stage072[202]}
   );
   gpc1_1 gpc1_1_2516(
      {stage072[69]},
      {stage072[203]}
   );
   gpc1_1 gpc1_1_2517(
      {stage072[70]},
      {stage072[204]}
   );
   gpc1_1 gpc1_1_2518(
      {stage072[71]},
      {stage072[205]}
   );
   gpc1_1 gpc1_1_2519(
      {stage072[72]},
      {stage072[206]}
   );
   gpc1_1 gpc1_1_2520(
      {stage072[73]},
      {stage072[207]}
   );
   gpc1_1 gpc1_1_2521(
      {stage072[74]},
      {stage072[208]}
   );
   gpc1_1 gpc1_1_2522(
      {stage072[75]},
      {stage072[209]}
   );
   gpc1_1 gpc1_1_2523(
      {stage072[76]},
      {stage072[210]}
   );
   gpc1_1 gpc1_1_2524(
      {stage072[77]},
      {stage072[211]}
   );
   gpc615_5 gpc615_5_2525(
      {stage072[78], stage072[79], stage072[80], stage072[81], stage072[82]},
      {stage073[18]},
      {stage074[0], stage074[1], stage074[2], stage074[3], stage074[4], stage074[5]},
      {stage076[128], stage075[131], stage074[136], stage073[150], stage072[212]}
   );
   gpc615_5 gpc615_5_2526(
      {stage072[83], stage072[84], stage072[85], stage072[86], stage072[87]},
      {stage073[19]},
      {stage074[6], stage074[7], stage074[8], stage074[9], stage074[10], stage074[11]},
      {stage076[129], stage075[132], stage074[137], stage073[151], stage072[213]}
   );
   gpc615_5 gpc615_5_2527(
      {stage072[88], stage072[89], stage072[90], stage072[91], stage072[92]},
      {stage073[20]},
      {stage074[12], stage074[13], stage074[14], stage074[15], stage074[16], stage074[17]},
      {stage076[130], stage075[133], stage074[138], stage073[152], stage072[214]}
   );
   gpc615_5 gpc615_5_2528(
      {stage072[93], stage072[94], stage072[95], stage072[96], stage072[97]},
      {stage073[21]},
      {stage074[18], stage074[19], stage074[20], stage074[21], stage074[22], stage074[23]},
      {stage076[131], stage075[134], stage074[139], stage073[153], stage072[215]}
   );
   gpc615_5 gpc615_5_2529(
      {stage072[98], stage072[99], stage072[100], stage072[101], stage072[102]},
      {stage073[22]},
      {stage074[24], stage074[25], stage074[26], stage074[27], stage074[28], stage074[29]},
      {stage076[132], stage075[135], stage074[140], stage073[154], stage072[216]}
   );
   gpc615_5 gpc615_5_2530(
      {stage072[103], stage072[104], stage072[105], stage072[106], stage072[107]},
      {stage073[23]},
      {stage074[30], stage074[31], stage074[32], stage074[33], stage074[34], stage074[35]},
      {stage076[133], stage075[136], stage074[141], stage073[155], stage072[217]}
   );
   gpc615_5 gpc615_5_2531(
      {stage072[108], stage072[109], stage072[110], stage072[111], stage072[112]},
      {stage073[24]},
      {stage074[36], stage074[37], stage074[38], stage074[39], stage074[40], stage074[41]},
      {stage076[134], stage075[137], stage074[142], stage073[156], stage072[218]}
   );
   gpc615_5 gpc615_5_2532(
      {stage072[113], stage072[114], stage072[115], stage072[116], stage072[117]},
      {stage073[25]},
      {stage074[42], stage074[43], stage074[44], stage074[45], stage074[46], stage074[47]},
      {stage076[135], stage075[138], stage074[143], stage073[157], stage072[219]}
   );
   gpc615_5 gpc615_5_2533(
      {stage072[118], stage072[119], stage072[120], stage072[121], stage072[122]},
      {stage073[26]},
      {stage074[48], stage074[49], stage074[50], stage074[51], stage074[52], stage074[53]},
      {stage076[136], stage075[139], stage074[144], stage073[158], stage072[220]}
   );
   gpc615_5 gpc615_5_2534(
      {stage072[123], stage072[124], stage072[125], stage072[126], stage072[127]},
      {stage073[27]},
      {stage074[54], stage074[55], stage074[56], stage074[57], stage074[58], stage074[59]},
      {stage076[137], stage075[140], stage074[145], stage073[159], stage072[221]}
   );
   gpc1_1 gpc1_1_2535(
      {stage073[28]},
      {stage073[160]}
   );
   gpc1_1 gpc1_1_2536(
      {stage073[29]},
      {stage073[161]}
   );
   gpc1_1 gpc1_1_2537(
      {stage073[30]},
      {stage073[162]}
   );
   gpc1_1 gpc1_1_2538(
      {stage073[31]},
      {stage073[163]}
   );
   gpc1_1 gpc1_1_2539(
      {stage073[32]},
      {stage073[164]}
   );
   gpc1_1 gpc1_1_2540(
      {stage073[33]},
      {stage073[165]}
   );
   gpc1_1 gpc1_1_2541(
      {stage073[34]},
      {stage073[166]}
   );
   gpc1_1 gpc1_1_2542(
      {stage073[35]},
      {stage073[167]}
   );
   gpc1_1 gpc1_1_2543(
      {stage073[36]},
      {stage073[168]}
   );
   gpc1_1 gpc1_1_2544(
      {stage073[37]},
      {stage073[169]}
   );
   gpc1_1 gpc1_1_2545(
      {stage073[38]},
      {stage073[170]}
   );
   gpc1_1 gpc1_1_2546(
      {stage073[39]},
      {stage073[171]}
   );
   gpc1_1 gpc1_1_2547(
      {stage073[40]},
      {stage073[172]}
   );
   gpc1_1 gpc1_1_2548(
      {stage073[41]},
      {stage073[173]}
   );
   gpc1_1 gpc1_1_2549(
      {stage073[42]},
      {stage073[174]}
   );
   gpc1_1 gpc1_1_2550(
      {stage073[43]},
      {stage073[175]}
   );
   gpc1_1 gpc1_1_2551(
      {stage073[44]},
      {stage073[176]}
   );
   gpc1_1 gpc1_1_2552(
      {stage073[45]},
      {stage073[177]}
   );
   gpc606_5 gpc606_5_2553(
      {stage073[46], stage073[47], stage073[48], stage073[49], stage073[50], stage073[51]},
      {stage075[0], stage075[1], stage075[2], stage075[3], stage075[4], stage075[5]},
      {stage077[128], stage076[138], stage075[141], stage074[146], stage073[178]}
   );
   gpc606_5 gpc606_5_2554(
      {stage073[52], stage073[53], stage073[54], stage073[55], stage073[56], stage073[57]},
      {stage075[6], stage075[7], stage075[8], stage075[9], stage075[10], stage075[11]},
      {stage077[129], stage076[139], stage075[142], stage074[147], stage073[179]}
   );
   gpc606_5 gpc606_5_2555(
      {stage073[58], stage073[59], stage073[60], stage073[61], stage073[62], stage073[63]},
      {stage075[12], stage075[13], stage075[14], stage075[15], stage075[16], stage075[17]},
      {stage077[130], stage076[140], stage075[143], stage074[148], stage073[180]}
   );
   gpc606_5 gpc606_5_2556(
      {stage073[64], stage073[65], stage073[66], stage073[67], stage073[68], stage073[69]},
      {stage075[18], stage075[19], stage075[20], stage075[21], stage075[22], stage075[23]},
      {stage077[131], stage076[141], stage075[144], stage074[149], stage073[181]}
   );
   gpc606_5 gpc606_5_2557(
      {stage073[70], stage073[71], stage073[72], stage073[73], stage073[74], stage073[75]},
      {stage075[24], stage075[25], stage075[26], stage075[27], stage075[28], stage075[29]},
      {stage077[132], stage076[142], stage075[145], stage074[150], stage073[182]}
   );
   gpc606_5 gpc606_5_2558(
      {stage073[76], stage073[77], stage073[78], stage073[79], stage073[80], stage073[81]},
      {stage075[30], stage075[31], stage075[32], stage075[33], stage075[34], stage075[35]},
      {stage077[133], stage076[143], stage075[146], stage074[151], stage073[183]}
   );
   gpc606_5 gpc606_5_2559(
      {stage073[82], stage073[83], stage073[84], stage073[85], stage073[86], stage073[87]},
      {stage075[36], stage075[37], stage075[38], stage075[39], stage075[40], stage075[41]},
      {stage077[134], stage076[144], stage075[147], stage074[152], stage073[184]}
   );
   gpc615_5 gpc615_5_2560(
      {stage073[88], stage073[89], stage073[90], stage073[91], stage073[92]},
      {stage074[60]},
      {stage075[42], stage075[43], stage075[44], stage075[45], stage075[46], stage075[47]},
      {stage077[135], stage076[145], stage075[148], stage074[153], stage073[185]}
   );
   gpc615_5 gpc615_5_2561(
      {stage073[93], stage073[94], stage073[95], stage073[96], stage073[97]},
      {stage074[61]},
      {stage075[48], stage075[49], stage075[50], stage075[51], stage075[52], stage075[53]},
      {stage077[136], stage076[146], stage075[149], stage074[154], stage073[186]}
   );
   gpc615_5 gpc615_5_2562(
      {stage073[98], stage073[99], stage073[100], stage073[101], stage073[102]},
      {stage074[62]},
      {stage075[54], stage075[55], stage075[56], stage075[57], stage075[58], stage075[59]},
      {stage077[137], stage076[147], stage075[150], stage074[155], stage073[187]}
   );
   gpc615_5 gpc615_5_2563(
      {stage073[103], stage073[104], stage073[105], stage073[106], stage073[107]},
      {stage074[63]},
      {stage075[60], stage075[61], stage075[62], stage075[63], stage075[64], stage075[65]},
      {stage077[138], stage076[148], stage075[151], stage074[156], stage073[188]}
   );
   gpc615_5 gpc615_5_2564(
      {stage073[108], stage073[109], stage073[110], stage073[111], stage073[112]},
      {stage074[64]},
      {stage075[66], stage075[67], stage075[68], stage075[69], stage075[70], stage075[71]},
      {stage077[139], stage076[149], stage075[152], stage074[157], stage073[189]}
   );
   gpc615_5 gpc615_5_2565(
      {stage073[113], stage073[114], stage073[115], stage073[116], stage073[117]},
      {stage074[65]},
      {stage075[72], stage075[73], stage075[74], stage075[75], stage075[76], stage075[77]},
      {stage077[140], stage076[150], stage075[153], stage074[158], stage073[190]}
   );
   gpc615_5 gpc615_5_2566(
      {stage073[118], stage073[119], stage073[120], stage073[121], stage073[122]},
      {stage074[66]},
      {stage075[78], stage075[79], stage075[80], stage075[81], stage075[82], stage075[83]},
      {stage077[141], stage076[151], stage075[154], stage074[159], stage073[191]}
   );
   gpc615_5 gpc615_5_2567(
      {stage073[123], stage073[124], stage073[125], stage073[126], stage073[127]},
      {stage074[67]},
      {stage075[84], stage075[85], stage075[86], stage075[87], stage075[88], stage075[89]},
      {stage077[142], stage076[152], stage075[155], stage074[160], stage073[192]}
   );
   gpc1_1 gpc1_1_2568(
      {stage074[68]},
      {stage074[161]}
   );
   gpc1_1 gpc1_1_2569(
      {stage074[69]},
      {stage074[162]}
   );
   gpc1_1 gpc1_1_2570(
      {stage074[70]},
      {stage074[163]}
   );
   gpc1_1 gpc1_1_2571(
      {stage074[71]},
      {stage074[164]}
   );
   gpc1_1 gpc1_1_2572(
      {stage074[72]},
      {stage074[165]}
   );
   gpc1_1 gpc1_1_2573(
      {stage074[73]},
      {stage074[166]}
   );
   gpc1_1 gpc1_1_2574(
      {stage074[74]},
      {stage074[167]}
   );
   gpc1_1 gpc1_1_2575(
      {stage074[75]},
      {stage074[168]}
   );
   gpc1_1 gpc1_1_2576(
      {stage074[76]},
      {stage074[169]}
   );
   gpc1_1 gpc1_1_2577(
      {stage074[77]},
      {stage074[170]}
   );
   gpc1_1 gpc1_1_2578(
      {stage074[78]},
      {stage074[171]}
   );
   gpc1_1 gpc1_1_2579(
      {stage074[79]},
      {stage074[172]}
   );
   gpc1_1 gpc1_1_2580(
      {stage074[80]},
      {stage074[173]}
   );
   gpc1_1 gpc1_1_2581(
      {stage074[81]},
      {stage074[174]}
   );
   gpc1_1 gpc1_1_2582(
      {stage074[82]},
      {stage074[175]}
   );
   gpc1_1 gpc1_1_2583(
      {stage074[83]},
      {stage074[176]}
   );
   gpc1_1 gpc1_1_2584(
      {stage074[84]},
      {stage074[177]}
   );
   gpc1_1 gpc1_1_2585(
      {stage074[85]},
      {stage074[178]}
   );
   gpc1_1 gpc1_1_2586(
      {stage074[86]},
      {stage074[179]}
   );
   gpc1_1 gpc1_1_2587(
      {stage074[87]},
      {stage074[180]}
   );
   gpc1_1 gpc1_1_2588(
      {stage074[88]},
      {stage074[181]}
   );
   gpc606_5 gpc606_5_2589(
      {stage074[89], stage074[90], stage074[91], stage074[92], stage074[93], stage074[94]},
      {stage076[0], stage076[1], stage076[2], stage076[3], stage076[4], stage076[5]},
      {stage078[128], stage077[143], stage076[153], stage075[156], stage074[182]}
   );
   gpc606_5 gpc606_5_2590(
      {stage074[95], stage074[96], stage074[97], stage074[98], stage074[99], stage074[100]},
      {stage076[6], stage076[7], stage076[8], stage076[9], stage076[10], stage076[11]},
      {stage078[129], stage077[144], stage076[154], stage075[157], stage074[183]}
   );
   gpc606_5 gpc606_5_2591(
      {stage074[101], stage074[102], stage074[103], stage074[104], stage074[105], stage074[106]},
      {stage076[12], stage076[13], stage076[14], stage076[15], stage076[16], stage076[17]},
      {stage078[130], stage077[145], stage076[155], stage075[158], stage074[184]}
   );
   gpc606_5 gpc606_5_2592(
      {stage074[107], stage074[108], stage074[109], stage074[110], stage074[111], stage074[112]},
      {stage076[18], stage076[19], stage076[20], stage076[21], stage076[22], stage076[23]},
      {stage078[131], stage077[146], stage076[156], stage075[159], stage074[185]}
   );
   gpc615_5 gpc615_5_2593(
      {stage074[113], stage074[114], stage074[115], stage074[116], stage074[117]},
      {stage075[90]},
      {stage076[24], stage076[25], stage076[26], stage076[27], stage076[28], stage076[29]},
      {stage078[132], stage077[147], stage076[157], stage075[160], stage074[186]}
   );
   gpc615_5 gpc615_5_2594(
      {stage074[118], stage074[119], stage074[120], stage074[121], stage074[122]},
      {stage075[91]},
      {stage076[30], stage076[31], stage076[32], stage076[33], stage076[34], stage076[35]},
      {stage078[133], stage077[148], stage076[158], stage075[161], stage074[187]}
   );
   gpc615_5 gpc615_5_2595(
      {stage074[123], stage074[124], stage074[125], stage074[126], stage074[127]},
      {stage075[92]},
      {stage076[36], stage076[37], stage076[38], stage076[39], stage076[40], stage076[41]},
      {stage078[134], stage077[149], stage076[159], stage075[162], stage074[188]}
   );
   gpc606_5 gpc606_5_2596(
      {stage075[93], stage075[94], stage075[95], stage075[96], stage075[97], stage075[98]},
      {stage077[0], stage077[1], stage077[2], stage077[3], stage077[4], stage077[5]},
      {stage079[128], stage078[135], stage077[150], stage076[160], stage075[163]}
   );
   gpc606_5 gpc606_5_2597(
      {stage075[99], stage075[100], stage075[101], stage075[102], stage075[103], stage075[104]},
      {stage077[6], stage077[7], stage077[8], stage077[9], stage077[10], stage077[11]},
      {stage079[129], stage078[136], stage077[151], stage076[161], stage075[164]}
   );
   gpc606_5 gpc606_5_2598(
      {stage075[105], stage075[106], stage075[107], stage075[108], stage075[109], stage075[110]},
      {stage077[12], stage077[13], stage077[14], stage077[15], stage077[16], stage077[17]},
      {stage079[130], stage078[137], stage077[152], stage076[162], stage075[165]}
   );
   gpc606_5 gpc606_5_2599(
      {stage075[111], stage075[112], stage075[113], stage075[114], stage075[115], stage075[116]},
      {stage077[18], stage077[19], stage077[20], stage077[21], stage077[22], stage077[23]},
      {stage079[131], stage078[138], stage077[153], stage076[163], stage075[166]}
   );
   gpc606_5 gpc606_5_2600(
      {stage075[117], stage075[118], stage075[119], stage075[120], stage075[121], stage075[122]},
      {stage077[24], stage077[25], stage077[26], stage077[27], stage077[28], stage077[29]},
      {stage079[132], stage078[139], stage077[154], stage076[164], stage075[167]}
   );
   gpc615_5 gpc615_5_2601(
      {stage075[123], stage075[124], stage075[125], stage075[126], stage075[127]},
      {stage076[42]},
      {stage077[30], stage077[31], stage077[32], stage077[33], stage077[34], stage077[35]},
      {stage079[133], stage078[140], stage077[155], stage076[165], stage075[168]}
   );
   gpc1_1 gpc1_1_2602(
      {stage076[43]},
      {stage076[166]}
   );
   gpc606_5 gpc606_5_2603(
      {stage076[44], stage076[45], stage076[46], stage076[47], stage076[48], stage076[49]},
      {stage078[0], stage078[1], stage078[2], stage078[3], stage078[4], stage078[5]},
      {stage080[128], stage079[134], stage078[141], stage077[156], stage076[167]}
   );
   gpc606_5 gpc606_5_2604(
      {stage076[50], stage076[51], stage076[52], stage076[53], stage076[54], stage076[55]},
      {stage078[6], stage078[7], stage078[8], stage078[9], stage078[10], stage078[11]},
      {stage080[129], stage079[135], stage078[142], stage077[157], stage076[168]}
   );
   gpc606_5 gpc606_5_2605(
      {stage076[56], stage076[57], stage076[58], stage076[59], stage076[60], stage076[61]},
      {stage078[12], stage078[13], stage078[14], stage078[15], stage078[16], stage078[17]},
      {stage080[130], stage079[136], stage078[143], stage077[158], stage076[169]}
   );
   gpc606_5 gpc606_5_2606(
      {stage076[62], stage076[63], stage076[64], stage076[65], stage076[66], stage076[67]},
      {stage078[18], stage078[19], stage078[20], stage078[21], stage078[22], stage078[23]},
      {stage080[131], stage079[137], stage078[144], stage077[159], stage076[170]}
   );
   gpc606_5 gpc606_5_2607(
      {stage076[68], stage076[69], stage076[70], stage076[71], stage076[72], stage076[73]},
      {stage078[24], stage078[25], stage078[26], stage078[27], stage078[28], stage078[29]},
      {stage080[132], stage079[138], stage078[145], stage077[160], stage076[171]}
   );
   gpc606_5 gpc606_5_2608(
      {stage076[74], stage076[75], stage076[76], stage076[77], stage076[78], stage076[79]},
      {stage078[30], stage078[31], stage078[32], stage078[33], stage078[34], stage078[35]},
      {stage080[133], stage079[139], stage078[146], stage077[161], stage076[172]}
   );
   gpc606_5 gpc606_5_2609(
      {stage076[80], stage076[81], stage076[82], stage076[83], stage076[84], stage076[85]},
      {stage078[36], stage078[37], stage078[38], stage078[39], stage078[40], stage078[41]},
      {stage080[134], stage079[140], stage078[147], stage077[162], stage076[173]}
   );
   gpc606_5 gpc606_5_2610(
      {stage076[86], stage076[87], stage076[88], stage076[89], stage076[90], stage076[91]},
      {stage078[42], stage078[43], stage078[44], stage078[45], stage078[46], stage078[47]},
      {stage080[135], stage079[141], stage078[148], stage077[163], stage076[174]}
   );
   gpc606_5 gpc606_5_2611(
      {stage076[92], stage076[93], stage076[94], stage076[95], stage076[96], stage076[97]},
      {stage078[48], stage078[49], stage078[50], stage078[51], stage078[52], stage078[53]},
      {stage080[136], stage079[142], stage078[149], stage077[164], stage076[175]}
   );
   gpc615_5 gpc615_5_2612(
      {stage076[98], stage076[99], stage076[100], stage076[101], stage076[102]},
      {stage077[36]},
      {stage078[54], stage078[55], stage078[56], stage078[57], stage078[58], stage078[59]},
      {stage080[137], stage079[143], stage078[150], stage077[165], stage076[176]}
   );
   gpc615_5 gpc615_5_2613(
      {stage076[103], stage076[104], stage076[105], stage076[106], stage076[107]},
      {stage077[37]},
      {stage078[60], stage078[61], stage078[62], stage078[63], stage078[64], stage078[65]},
      {stage080[138], stage079[144], stage078[151], stage077[166], stage076[177]}
   );
   gpc615_5 gpc615_5_2614(
      {stage076[108], stage076[109], stage076[110], stage076[111], stage076[112]},
      {stage077[38]},
      {stage078[66], stage078[67], stage078[68], stage078[69], stage078[70], stage078[71]},
      {stage080[139], stage079[145], stage078[152], stage077[167], stage076[178]}
   );
   gpc615_5 gpc615_5_2615(
      {stage076[113], stage076[114], stage076[115], stage076[116], stage076[117]},
      {stage077[39]},
      {stage078[72], stage078[73], stage078[74], stage078[75], stage078[76], stage078[77]},
      {stage080[140], stage079[146], stage078[153], stage077[168], stage076[179]}
   );
   gpc615_5 gpc615_5_2616(
      {stage076[118], stage076[119], stage076[120], stage076[121], stage076[122]},
      {stage077[40]},
      {stage078[78], stage078[79], stage078[80], stage078[81], stage078[82], stage078[83]},
      {stage080[141], stage079[147], stage078[154], stage077[169], stage076[180]}
   );
   gpc615_5 gpc615_5_2617(
      {stage076[123], stage076[124], stage076[125], stage076[126], stage076[127]},
      {stage077[41]},
      {stage078[84], stage078[85], stage078[86], stage078[87], stage078[88], stage078[89]},
      {stage080[142], stage079[148], stage078[155], stage077[170], stage076[181]}
   );
   gpc1_1 gpc1_1_2618(
      {stage077[42]},
      {stage077[171]}
   );
   gpc1_1 gpc1_1_2619(
      {stage077[43]},
      {stage077[172]}
   );
   gpc1_1 gpc1_1_2620(
      {stage077[44]},
      {stage077[173]}
   );
   gpc1_1 gpc1_1_2621(
      {stage077[45]},
      {stage077[174]}
   );
   gpc1_1 gpc1_1_2622(
      {stage077[46]},
      {stage077[175]}
   );
   gpc1_1 gpc1_1_2623(
      {stage077[47]},
      {stage077[176]}
   );
   gpc1_1 gpc1_1_2624(
      {stage077[48]},
      {stage077[177]}
   );
   gpc1_1 gpc1_1_2625(
      {stage077[49]},
      {stage077[178]}
   );
   gpc1_1 gpc1_1_2626(
      {stage077[50]},
      {stage077[179]}
   );
   gpc1_1 gpc1_1_2627(
      {stage077[51]},
      {stage077[180]}
   );
   gpc1_1 gpc1_1_2628(
      {stage077[52]},
      {stage077[181]}
   );
   gpc1_1 gpc1_1_2629(
      {stage077[53]},
      {stage077[182]}
   );
   gpc1_1 gpc1_1_2630(
      {stage077[54]},
      {stage077[183]}
   );
   gpc1_1 gpc1_1_2631(
      {stage077[55]},
      {stage077[184]}
   );
   gpc1_1 gpc1_1_2632(
      {stage077[56]},
      {stage077[185]}
   );
   gpc1_1 gpc1_1_2633(
      {stage077[57]},
      {stage077[186]}
   );
   gpc1_1 gpc1_1_2634(
      {stage077[58]},
      {stage077[187]}
   );
   gpc1_1 gpc1_1_2635(
      {stage077[59]},
      {stage077[188]}
   );
   gpc1_1 gpc1_1_2636(
      {stage077[60]},
      {stage077[189]}
   );
   gpc1_1 gpc1_1_2637(
      {stage077[61]},
      {stage077[190]}
   );
   gpc1_1 gpc1_1_2638(
      {stage077[62]},
      {stage077[191]}
   );
   gpc7_3 gpc7_3_2639(
      {stage077[63], stage077[64], stage077[65], stage077[66], stage077[67], stage077[68], stage077[69]},
      {stage079[149], stage078[156], stage077[192]}
   );
   gpc7_3 gpc7_3_2640(
      {stage077[70], stage077[71], stage077[72], stage077[73], stage077[74], stage077[75], stage077[76]},
      {stage079[150], stage078[157], stage077[193]}
   );
   gpc606_5 gpc606_5_2641(
      {stage077[77], stage077[78], stage077[79], stage077[80], stage077[81], stage077[82]},
      {stage079[0], stage079[1], stage079[2], stage079[3], stage079[4], stage079[5]},
      {stage081[128], stage080[143], stage079[151], stage078[158], stage077[194]}
   );
   gpc606_5 gpc606_5_2642(
      {stage077[83], stage077[84], stage077[85], stage077[86], stage077[87], stage077[88]},
      {stage079[6], stage079[7], stage079[8], stage079[9], stage079[10], stage079[11]},
      {stage081[129], stage080[144], stage079[152], stage078[159], stage077[195]}
   );
   gpc606_5 gpc606_5_2643(
      {stage077[89], stage077[90], stage077[91], stage077[92], stage077[93], stage077[94]},
      {stage079[12], stage079[13], stage079[14], stage079[15], stage079[16], stage079[17]},
      {stage081[130], stage080[145], stage079[153], stage078[160], stage077[196]}
   );
   gpc606_5 gpc606_5_2644(
      {stage077[95], stage077[96], stage077[97], stage077[98], stage077[99], stage077[100]},
      {stage079[18], stage079[19], stage079[20], stage079[21], stage079[22], stage079[23]},
      {stage081[131], stage080[146], stage079[154], stage078[161], stage077[197]}
   );
   gpc606_5 gpc606_5_2645(
      {stage077[101], stage077[102], stage077[103], stage077[104], stage077[105], stage077[106]},
      {stage079[24], stage079[25], stage079[26], stage079[27], stage079[28], stage079[29]},
      {stage081[132], stage080[147], stage079[155], stage078[162], stage077[198]}
   );
   gpc606_5 gpc606_5_2646(
      {stage077[107], stage077[108], stage077[109], stage077[110], stage077[111], stage077[112]},
      {stage079[30], stage079[31], stage079[32], stage079[33], stage079[34], stage079[35]},
      {stage081[133], stage080[148], stage079[156], stage078[163], stage077[199]}
   );
   gpc615_5 gpc615_5_2647(
      {stage077[113], stage077[114], stage077[115], stage077[116], stage077[117]},
      {stage078[90]},
      {stage079[36], stage079[37], stage079[38], stage079[39], stage079[40], stage079[41]},
      {stage081[134], stage080[149], stage079[157], stage078[164], stage077[200]}
   );
   gpc615_5 gpc615_5_2648(
      {stage077[118], stage077[119], stage077[120], stage077[121], stage077[122]},
      {stage078[91]},
      {stage079[42], stage079[43], stage079[44], stage079[45], stage079[46], stage079[47]},
      {stage081[135], stage080[150], stage079[158], stage078[165], stage077[201]}
   );
   gpc615_5 gpc615_5_2649(
      {stage077[123], stage077[124], stage077[125], stage077[126], stage077[127]},
      {stage078[92]},
      {stage079[48], stage079[49], stage079[50], stage079[51], stage079[52], stage079[53]},
      {stage081[136], stage080[151], stage079[159], stage078[166], stage077[202]}
   );
   gpc606_5 gpc606_5_2650(
      {stage078[93], stage078[94], stage078[95], stage078[96], stage078[97], stage078[98]},
      {stage080[0], stage080[1], stage080[2], stage080[3], stage080[4], stage080[5]},
      {stage082[128], stage081[137], stage080[152], stage079[160], stage078[167]}
   );
   gpc615_5 gpc615_5_2651(
      {stage078[99], stage078[100], stage078[101], stage078[102], stage078[103]},
      {stage079[54]},
      {stage080[6], stage080[7], stage080[8], stage080[9], stage080[10], stage080[11]},
      {stage082[129], stage081[138], stage080[153], stage079[161], stage078[168]}
   );
   gpc615_5 gpc615_5_2652(
      {stage078[104], stage078[105], stage078[106], stage078[107], stage078[108]},
      {stage079[55]},
      {stage080[12], stage080[13], stage080[14], stage080[15], stage080[16], stage080[17]},
      {stage082[130], stage081[139], stage080[154], stage079[162], stage078[169]}
   );
   gpc615_5 gpc615_5_2653(
      {stage078[109], stage078[110], stage078[111], stage078[112], stage078[113]},
      {stage079[56]},
      {stage080[18], stage080[19], stage080[20], stage080[21], stage080[22], stage080[23]},
      {stage082[131], stage081[140], stage080[155], stage079[163], stage078[170]}
   );
   gpc615_5 gpc615_5_2654(
      {stage078[114], stage078[115], stage078[116], stage078[117], stage078[118]},
      {stage079[57]},
      {stage080[24], stage080[25], stage080[26], stage080[27], stage080[28], stage080[29]},
      {stage082[132], stage081[141], stage080[156], stage079[164], stage078[171]}
   );
   gpc615_5 gpc615_5_2655(
      {stage078[119], stage078[120], stage078[121], stage078[122], stage078[123]},
      {stage079[58]},
      {stage080[30], stage080[31], stage080[32], stage080[33], stage080[34], stage080[35]},
      {stage082[133], stage081[142], stage080[157], stage079[165], stage078[172]}
   );
   gpc615_5 gpc615_5_2656(
      {stage078[124], stage078[125], stage078[126], stage078[127], 1'h0},
      {stage079[59]},
      {stage080[36], stage080[37], stage080[38], stage080[39], stage080[40], stage080[41]},
      {stage082[134], stage081[143], stage080[158], stage079[166], stage078[173]}
   );
   gpc1_1 gpc1_1_2657(
      {stage079[60]},
      {stage079[167]}
   );
   gpc1_1 gpc1_1_2658(
      {stage079[61]},
      {stage079[168]}
   );
   gpc1_1 gpc1_1_2659(
      {stage079[62]},
      {stage079[169]}
   );
   gpc1_1 gpc1_1_2660(
      {stage079[63]},
      {stage079[170]}
   );
   gpc1_1 gpc1_1_2661(
      {stage079[64]},
      {stage079[171]}
   );
   gpc1_1 gpc1_1_2662(
      {stage079[65]},
      {stage079[172]}
   );
   gpc615_5 gpc615_5_2663(
      {stage079[66], stage079[67], stage079[68], stage079[69], stage079[70]},
      {stage080[42]},
      {stage081[0], stage081[1], stage081[2], stage081[3], stage081[4], stage081[5]},
      {stage083[128], stage082[135], stage081[144], stage080[159], stage079[173]}
   );
   gpc615_5 gpc615_5_2664(
      {stage079[71], stage079[72], stage079[73], stage079[74], stage079[75]},
      {stage080[43]},
      {stage081[6], stage081[7], stage081[8], stage081[9], stage081[10], stage081[11]},
      {stage083[129], stage082[136], stage081[145], stage080[160], stage079[174]}
   );
   gpc615_5 gpc615_5_2665(
      {stage079[76], stage079[77], stage079[78], stage079[79], stage079[80]},
      {stage080[44]},
      {stage081[12], stage081[13], stage081[14], stage081[15], stage081[16], stage081[17]},
      {stage083[130], stage082[137], stage081[146], stage080[161], stage079[175]}
   );
   gpc615_5 gpc615_5_2666(
      {stage079[81], stage079[82], stage079[83], stage079[84], stage079[85]},
      {stage080[45]},
      {stage081[18], stage081[19], stage081[20], stage081[21], stage081[22], stage081[23]},
      {stage083[131], stage082[138], stage081[147], stage080[162], stage079[176]}
   );
   gpc615_5 gpc615_5_2667(
      {stage079[86], stage079[87], stage079[88], stage079[89], stage079[90]},
      {stage080[46]},
      {stage081[24], stage081[25], stage081[26], stage081[27], stage081[28], stage081[29]},
      {stage083[132], stage082[139], stage081[148], stage080[163], stage079[177]}
   );
   gpc615_5 gpc615_5_2668(
      {stage079[91], stage079[92], stage079[93], stage079[94], stage079[95]},
      {stage080[47]},
      {stage081[30], stage081[31], stage081[32], stage081[33], stage081[34], stage081[35]},
      {stage083[133], stage082[140], stage081[149], stage080[164], stage079[178]}
   );
   gpc615_5 gpc615_5_2669(
      {stage079[96], stage079[97], stage079[98], stage079[99], stage079[100]},
      {stage080[48]},
      {stage081[36], stage081[37], stage081[38], stage081[39], stage081[40], stage081[41]},
      {stage083[134], stage082[141], stage081[150], stage080[165], stage079[179]}
   );
   gpc615_5 gpc615_5_2670(
      {stage079[101], stage079[102], stage079[103], stage079[104], stage079[105]},
      {stage080[49]},
      {stage081[42], stage081[43], stage081[44], stage081[45], stage081[46], stage081[47]},
      {stage083[135], stage082[142], stage081[151], stage080[166], stage079[180]}
   );
   gpc615_5 gpc615_5_2671(
      {stage079[106], stage079[107], stage079[108], stage079[109], stage079[110]},
      {stage080[50]},
      {stage081[48], stage081[49], stage081[50], stage081[51], stage081[52], stage081[53]},
      {stage083[136], stage082[143], stage081[152], stage080[167], stage079[181]}
   );
   gpc615_5 gpc615_5_2672(
      {stage079[111], stage079[112], stage079[113], stage079[114], stage079[115]},
      {stage080[51]},
      {stage081[54], stage081[55], stage081[56], stage081[57], stage081[58], stage081[59]},
      {stage083[137], stage082[144], stage081[153], stage080[168], stage079[182]}
   );
   gpc1343_5 gpc1343_5_2673(
      {stage079[116], stage079[117], stage079[118]},
      {stage080[52], stage080[53], stage080[54], stage080[55]},
      {stage081[60], stage081[61], stage081[62]},
      {stage082[0]},
      {stage083[138], stage082[145], stage081[154], stage080[169], stage079[183]}
   );
   gpc1343_5 gpc1343_5_2674(
      {stage079[119], stage079[120], stage079[121]},
      {stage080[56], stage080[57], stage080[58], stage080[59]},
      {stage081[63], stage081[64], stage081[65]},
      {stage082[1]},
      {stage083[139], stage082[146], stage081[155], stage080[170], stage079[184]}
   );
   gpc1343_5 gpc1343_5_2675(
      {stage079[122], stage079[123], stage079[124]},
      {stage080[60], stage080[61], stage080[62], stage080[63]},
      {stage081[66], stage081[67], stage081[68]},
      {stage082[2]},
      {stage083[140], stage082[147], stage081[156], stage080[171], stage079[185]}
   );
   gpc1343_5 gpc1343_5_2676(
      {stage079[125], stage079[126], stage079[127]},
      {stage080[64], stage080[65], stage080[66], stage080[67]},
      {stage081[69], stage081[70], stage081[71]},
      {stage082[3]},
      {stage083[141], stage082[148], stage081[157], stage080[172], stage079[186]}
   );
   gpc1_1 gpc1_1_2677(
      {stage080[68]},
      {stage080[173]}
   );
   gpc1_1 gpc1_1_2678(
      {stage080[69]},
      {stage080[174]}
   );
   gpc1_1 gpc1_1_2679(
      {stage080[70]},
      {stage080[175]}
   );
   gpc1_1 gpc1_1_2680(
      {stage080[71]},
      {stage080[176]}
   );
   gpc1_1 gpc1_1_2681(
      {stage080[72]},
      {stage080[177]}
   );
   gpc1_1 gpc1_1_2682(
      {stage080[73]},
      {stage080[178]}
   );
   gpc1_1 gpc1_1_2683(
      {stage080[74]},
      {stage080[179]}
   );
   gpc1_1 gpc1_1_2684(
      {stage080[75]},
      {stage080[180]}
   );
   gpc1_1 gpc1_1_2685(
      {stage080[76]},
      {stage080[181]}
   );
   gpc1_1 gpc1_1_2686(
      {stage080[77]},
      {stage080[182]}
   );
   gpc1_1 gpc1_1_2687(
      {stage080[78]},
      {stage080[183]}
   );
   gpc1_1 gpc1_1_2688(
      {stage080[79]},
      {stage080[184]}
   );
   gpc1_1 gpc1_1_2689(
      {stage080[80]},
      {stage080[185]}
   );
   gpc1_1 gpc1_1_2690(
      {stage080[81]},
      {stage080[186]}
   );
   gpc1_1 gpc1_1_2691(
      {stage080[82]},
      {stage080[187]}
   );
   gpc1_1 gpc1_1_2692(
      {stage080[83]},
      {stage080[188]}
   );
   gpc1_1 gpc1_1_2693(
      {stage080[84]},
      {stage080[189]}
   );
   gpc1_1 gpc1_1_2694(
      {stage080[85]},
      {stage080[190]}
   );
   gpc1_1 gpc1_1_2695(
      {stage080[86]},
      {stage080[191]}
   );
   gpc1_1 gpc1_1_2696(
      {stage080[87]},
      {stage080[192]}
   );
   gpc1_1 gpc1_1_2697(
      {stage080[88]},
      {stage080[193]}
   );
   gpc1_1 gpc1_1_2698(
      {stage080[89]},
      {stage080[194]}
   );
   gpc1_1 gpc1_1_2699(
      {stage080[90]},
      {stage080[195]}
   );
   gpc606_5 gpc606_5_2700(
      {stage080[91], stage080[92], stage080[93], stage080[94], stage080[95], stage080[96]},
      {stage082[4], stage082[5], stage082[6], stage082[7], stage082[8], stage082[9]},
      {stage084[128], stage083[142], stage082[149], stage081[158], stage080[196]}
   );
   gpc606_5 gpc606_5_2701(
      {stage080[97], stage080[98], stage080[99], stage080[100], stage080[101], stage080[102]},
      {stage082[10], stage082[11], stage082[12], stage082[13], stage082[14], stage082[15]},
      {stage084[129], stage083[143], stage082[150], stage081[159], stage080[197]}
   );
   gpc615_5 gpc615_5_2702(
      {stage080[103], stage080[104], stage080[105], stage080[106], stage080[107]},
      {stage081[72]},
      {stage082[16], stage082[17], stage082[18], stage082[19], stage082[20], stage082[21]},
      {stage084[130], stage083[144], stage082[151], stage081[160], stage080[198]}
   );
   gpc615_5 gpc615_5_2703(
      {stage080[108], stage080[109], stage080[110], stage080[111], stage080[112]},
      {stage081[73]},
      {stage082[22], stage082[23], stage082[24], stage082[25], stage082[26], stage082[27]},
      {stage084[131], stage083[145], stage082[152], stage081[161], stage080[199]}
   );
   gpc615_5 gpc615_5_2704(
      {stage080[113], stage080[114], stage080[115], stage080[116], stage080[117]},
      {stage081[74]},
      {stage082[28], stage082[29], stage082[30], stage082[31], stage082[32], stage082[33]},
      {stage084[132], stage083[146], stage082[153], stage081[162], stage080[200]}
   );
   gpc615_5 gpc615_5_2705(
      {stage080[118], stage080[119], stage080[120], stage080[121], stage080[122]},
      {stage081[75]},
      {stage082[34], stage082[35], stage082[36], stage082[37], stage082[38], stage082[39]},
      {stage084[133], stage083[147], stage082[154], stage081[163], stage080[201]}
   );
   gpc615_5 gpc615_5_2706(
      {stage080[123], stage080[124], stage080[125], stage080[126], stage080[127]},
      {stage081[76]},
      {stage082[40], stage082[41], stage082[42], stage082[43], stage082[44], stage082[45]},
      {stage084[134], stage083[148], stage082[155], stage081[164], stage080[202]}
   );
   gpc1_1 gpc1_1_2707(
      {stage081[77]},
      {stage081[165]}
   );
   gpc606_5 gpc606_5_2708(
      {stage081[78], stage081[79], stage081[80], stage081[81], stage081[82], stage081[83]},
      {stage083[0], stage083[1], stage083[2], stage083[3], stage083[4], stage083[5]},
      {stage085[128], stage084[135], stage083[149], stage082[156], stage081[166]}
   );
   gpc606_5 gpc606_5_2709(
      {stage081[84], stage081[85], stage081[86], stage081[87], stage081[88], stage081[89]},
      {stage083[6], stage083[7], stage083[8], stage083[9], stage083[10], stage083[11]},
      {stage085[129], stage084[136], stage083[150], stage082[157], stage081[167]}
   );
   gpc606_5 gpc606_5_2710(
      {stage081[90], stage081[91], stage081[92], stage081[93], stage081[94], stage081[95]},
      {stage083[12], stage083[13], stage083[14], stage083[15], stage083[16], stage083[17]},
      {stage085[130], stage084[137], stage083[151], stage082[158], stage081[168]}
   );
   gpc606_5 gpc606_5_2711(
      {stage081[96], stage081[97], stage081[98], stage081[99], stage081[100], stage081[101]},
      {stage083[18], stage083[19], stage083[20], stage083[21], stage083[22], stage083[23]},
      {stage085[131], stage084[138], stage083[152], stage082[159], stage081[169]}
   );
   gpc606_5 gpc606_5_2712(
      {stage081[102], stage081[103], stage081[104], stage081[105], stage081[106], stage081[107]},
      {stage083[24], stage083[25], stage083[26], stage083[27], stage083[28], stage083[29]},
      {stage085[132], stage084[139], stage083[153], stage082[160], stage081[170]}
   );
   gpc615_5 gpc615_5_2713(
      {stage081[108], stage081[109], stage081[110], stage081[111], stage081[112]},
      {stage082[46]},
      {stage083[30], stage083[31], stage083[32], stage083[33], stage083[34], stage083[35]},
      {stage085[133], stage084[140], stage083[154], stage082[161], stage081[171]}
   );
   gpc615_5 gpc615_5_2714(
      {stage081[113], stage081[114], stage081[115], stage081[116], stage081[117]},
      {stage082[47]},
      {stage083[36], stage083[37], stage083[38], stage083[39], stage083[40], stage083[41]},
      {stage085[134], stage084[141], stage083[155], stage082[162], stage081[172]}
   );
   gpc615_5 gpc615_5_2715(
      {stage081[118], stage081[119], stage081[120], stage081[121], stage081[122]},
      {stage082[48]},
      {stage083[42], stage083[43], stage083[44], stage083[45], stage083[46], stage083[47]},
      {stage085[135], stage084[142], stage083[156], stage082[163], stage081[173]}
   );
   gpc615_5 gpc615_5_2716(
      {stage081[123], stage081[124], stage081[125], stage081[126], stage081[127]},
      {stage082[49]},
      {stage083[48], stage083[49], stage083[50], stage083[51], stage083[52], stage083[53]},
      {stage085[136], stage084[143], stage083[157], stage082[164], stage081[174]}
   );
   gpc1_1 gpc1_1_2717(
      {stage082[50]},
      {stage082[165]}
   );
   gpc1_1 gpc1_1_2718(
      {stage082[51]},
      {stage082[166]}
   );
   gpc1_1 gpc1_1_2719(
      {stage082[52]},
      {stage082[167]}
   );
   gpc1_1 gpc1_1_2720(
      {stage082[53]},
      {stage082[168]}
   );
   gpc1_1 gpc1_1_2721(
      {stage082[54]},
      {stage082[169]}
   );
   gpc1_1 gpc1_1_2722(
      {stage082[55]},
      {stage082[170]}
   );
   gpc1_1 gpc1_1_2723(
      {stage082[56]},
      {stage082[171]}
   );
   gpc1_1 gpc1_1_2724(
      {stage082[57]},
      {stage082[172]}
   );
   gpc1_1 gpc1_1_2725(
      {stage082[58]},
      {stage082[173]}
   );
   gpc1_1 gpc1_1_2726(
      {stage082[59]},
      {stage082[174]}
   );
   gpc1_1 gpc1_1_2727(
      {stage082[60]},
      {stage082[175]}
   );
   gpc1_1 gpc1_1_2728(
      {stage082[61]},
      {stage082[176]}
   );
   gpc1_1 gpc1_1_2729(
      {stage082[62]},
      {stage082[177]}
   );
   gpc1_1 gpc1_1_2730(
      {stage082[63]},
      {stage082[178]}
   );
   gpc1_1 gpc1_1_2731(
      {stage082[64]},
      {stage082[179]}
   );
   gpc1_1 gpc1_1_2732(
      {stage082[65]},
      {stage082[180]}
   );
   gpc1_1 gpc1_1_2733(
      {stage082[66]},
      {stage082[181]}
   );
   gpc1_1 gpc1_1_2734(
      {stage082[67]},
      {stage082[182]}
   );
   gpc1_1 gpc1_1_2735(
      {stage082[68]},
      {stage082[183]}
   );
   gpc1_1 gpc1_1_2736(
      {stage082[69]},
      {stage082[184]}
   );
   gpc1_1 gpc1_1_2737(
      {stage082[70]},
      {stage082[185]}
   );
   gpc1_1 gpc1_1_2738(
      {stage082[71]},
      {stage082[186]}
   );
   gpc1_1 gpc1_1_2739(
      {stage082[72]},
      {stage082[187]}
   );
   gpc1_1 gpc1_1_2740(
      {stage082[73]},
      {stage082[188]}
   );
   gpc1_1 gpc1_1_2741(
      {stage082[74]},
      {stage082[189]}
   );
   gpc1_1 gpc1_1_2742(
      {stage082[75]},
      {stage082[190]}
   );
   gpc1_1 gpc1_1_2743(
      {stage082[76]},
      {stage082[191]}
   );
   gpc1_1 gpc1_1_2744(
      {stage082[77]},
      {stage082[192]}
   );
   gpc1_1 gpc1_1_2745(
      {stage082[78]},
      {stage082[193]}
   );
   gpc1_1 gpc1_1_2746(
      {stage082[79]},
      {stage082[194]}
   );
   gpc1_1 gpc1_1_2747(
      {stage082[80]},
      {stage082[195]}
   );
   gpc1_1 gpc1_1_2748(
      {stage082[81]},
      {stage082[196]}
   );
   gpc1_1 gpc1_1_2749(
      {stage082[82]},
      {stage082[197]}
   );
   gpc1_1 gpc1_1_2750(
      {stage082[83]},
      {stage082[198]}
   );
   gpc1_1 gpc1_1_2751(
      {stage082[84]},
      {stage082[199]}
   );
   gpc1_1 gpc1_1_2752(
      {stage082[85]},
      {stage082[200]}
   );
   gpc1_1 gpc1_1_2753(
      {stage082[86]},
      {stage082[201]}
   );
   gpc1_1 gpc1_1_2754(
      {stage082[87]},
      {stage082[202]}
   );
   gpc1_1 gpc1_1_2755(
      {stage082[88]},
      {stage082[203]}
   );
   gpc1_1 gpc1_1_2756(
      {stage082[89]},
      {stage082[204]}
   );
   gpc1_1 gpc1_1_2757(
      {stage082[90]},
      {stage082[205]}
   );
   gpc1_1 gpc1_1_2758(
      {stage082[91]},
      {stage082[206]}
   );
   gpc1_1 gpc1_1_2759(
      {stage082[92]},
      {stage082[207]}
   );
   gpc615_5 gpc615_5_2760(
      {stage082[93], stage082[94], stage082[95], stage082[96], stage082[97]},
      {stage083[54]},
      {stage084[0], stage084[1], stage084[2], stage084[3], stage084[4], stage084[5]},
      {stage086[128], stage085[137], stage084[144], stage083[158], stage082[208]}
   );
   gpc615_5 gpc615_5_2761(
      {stage082[98], stage082[99], stage082[100], stage082[101], stage082[102]},
      {stage083[55]},
      {stage084[6], stage084[7], stage084[8], stage084[9], stage084[10], stage084[11]},
      {stage086[129], stage085[138], stage084[145], stage083[159], stage082[209]}
   );
   gpc615_5 gpc615_5_2762(
      {stage082[103], stage082[104], stage082[105], stage082[106], stage082[107]},
      {stage083[56]},
      {stage084[12], stage084[13], stage084[14], stage084[15], stage084[16], stage084[17]},
      {stage086[130], stage085[139], stage084[146], stage083[160], stage082[210]}
   );
   gpc615_5 gpc615_5_2763(
      {stage082[108], stage082[109], stage082[110], stage082[111], stage082[112]},
      {stage083[57]},
      {stage084[18], stage084[19], stage084[20], stage084[21], stage084[22], stage084[23]},
      {stage086[131], stage085[140], stage084[147], stage083[161], stage082[211]}
   );
   gpc615_5 gpc615_5_2764(
      {stage082[113], stage082[114], stage082[115], stage082[116], stage082[117]},
      {stage083[58]},
      {stage084[24], stage084[25], stage084[26], stage084[27], stage084[28], stage084[29]},
      {stage086[132], stage085[141], stage084[148], stage083[162], stage082[212]}
   );
   gpc615_5 gpc615_5_2765(
      {stage082[118], stage082[119], stage082[120], stage082[121], stage082[122]},
      {stage083[59]},
      {stage084[30], stage084[31], stage084[32], stage084[33], stage084[34], stage084[35]},
      {stage086[133], stage085[142], stage084[149], stage083[163], stage082[213]}
   );
   gpc615_5 gpc615_5_2766(
      {stage082[123], stage082[124], stage082[125], stage082[126], stage082[127]},
      {stage083[60]},
      {stage084[36], stage084[37], stage084[38], stage084[39], stage084[40], stage084[41]},
      {stage086[134], stage085[143], stage084[150], stage083[164], stage082[214]}
   );
   gpc1_1 gpc1_1_2767(
      {stage083[61]},
      {stage083[165]}
   );
   gpc1_1 gpc1_1_2768(
      {stage083[62]},
      {stage083[166]}
   );
   gpc1_1 gpc1_1_2769(
      {stage083[63]},
      {stage083[167]}
   );
   gpc1_1 gpc1_1_2770(
      {stage083[64]},
      {stage083[168]}
   );
   gpc1_1 gpc1_1_2771(
      {stage083[65]},
      {stage083[169]}
   );
   gpc1_1 gpc1_1_2772(
      {stage083[66]},
      {stage083[170]}
   );
   gpc1_1 gpc1_1_2773(
      {stage083[67]},
      {stage083[171]}
   );
   gpc1_1 gpc1_1_2774(
      {stage083[68]},
      {stage083[172]}
   );
   gpc1_1 gpc1_1_2775(
      {stage083[69]},
      {stage083[173]}
   );
   gpc1_1 gpc1_1_2776(
      {stage083[70]},
      {stage083[174]}
   );
   gpc1_1 gpc1_1_2777(
      {stage083[71]},
      {stage083[175]}
   );
   gpc1_1 gpc1_1_2778(
      {stage083[72]},
      {stage083[176]}
   );
   gpc1_1 gpc1_1_2779(
      {stage083[73]},
      {stage083[177]}
   );
   gpc1_1 gpc1_1_2780(
      {stage083[74]},
      {stage083[178]}
   );
   gpc1_1 gpc1_1_2781(
      {stage083[75]},
      {stage083[179]}
   );
   gpc1_1 gpc1_1_2782(
      {stage083[76]},
      {stage083[180]}
   );
   gpc1_1 gpc1_1_2783(
      {stage083[77]},
      {stage083[181]}
   );
   gpc1_1 gpc1_1_2784(
      {stage083[78]},
      {stage083[182]}
   );
   gpc1_1 gpc1_1_2785(
      {stage083[79]},
      {stage083[183]}
   );
   gpc1_1 gpc1_1_2786(
      {stage083[80]},
      {stage083[184]}
   );
   gpc1_1 gpc1_1_2787(
      {stage083[81]},
      {stage083[185]}
   );
   gpc1_1 gpc1_1_2788(
      {stage083[82]},
      {stage083[186]}
   );
   gpc615_5 gpc615_5_2789(
      {stage083[83], stage083[84], stage083[85], stage083[86], stage083[87]},
      {stage084[42]},
      {stage085[0], stage085[1], stage085[2], stage085[3], stage085[4], stage085[5]},
      {stage087[128], stage086[135], stage085[144], stage084[151], stage083[187]}
   );
   gpc615_5 gpc615_5_2790(
      {stage083[88], stage083[89], stage083[90], stage083[91], stage083[92]},
      {stage084[43]},
      {stage085[6], stage085[7], stage085[8], stage085[9], stage085[10], stage085[11]},
      {stage087[129], stage086[136], stage085[145], stage084[152], stage083[188]}
   );
   gpc615_5 gpc615_5_2791(
      {stage083[93], stage083[94], stage083[95], stage083[96], stage083[97]},
      {stage084[44]},
      {stage085[12], stage085[13], stage085[14], stage085[15], stage085[16], stage085[17]},
      {stage087[130], stage086[137], stage085[146], stage084[153], stage083[189]}
   );
   gpc615_5 gpc615_5_2792(
      {stage083[98], stage083[99], stage083[100], stage083[101], stage083[102]},
      {stage084[45]},
      {stage085[18], stage085[19], stage085[20], stage085[21], stage085[22], stage085[23]},
      {stage087[131], stage086[138], stage085[147], stage084[154], stage083[190]}
   );
   gpc615_5 gpc615_5_2793(
      {stage083[103], stage083[104], stage083[105], stage083[106], stage083[107]},
      {stage084[46]},
      {stage085[24], stage085[25], stage085[26], stage085[27], stage085[28], stage085[29]},
      {stage087[132], stage086[139], stage085[148], stage084[155], stage083[191]}
   );
   gpc615_5 gpc615_5_2794(
      {stage083[108], stage083[109], stage083[110], stage083[111], stage083[112]},
      {stage084[47]},
      {stage085[30], stage085[31], stage085[32], stage085[33], stage085[34], stage085[35]},
      {stage087[133], stage086[140], stage085[149], stage084[156], stage083[192]}
   );
   gpc615_5 gpc615_5_2795(
      {stage083[113], stage083[114], stage083[115], stage083[116], stage083[117]},
      {stage084[48]},
      {stage085[36], stage085[37], stage085[38], stage085[39], stage085[40], stage085[41]},
      {stage087[134], stage086[141], stage085[150], stage084[157], stage083[193]}
   );
   gpc615_5 gpc615_5_2796(
      {stage083[118], stage083[119], stage083[120], stage083[121], stage083[122]},
      {stage084[49]},
      {stage085[42], stage085[43], stage085[44], stage085[45], stage085[46], stage085[47]},
      {stage087[135], stage086[142], stage085[151], stage084[158], stage083[194]}
   );
   gpc615_5 gpc615_5_2797(
      {stage083[123], stage083[124], stage083[125], stage083[126], stage083[127]},
      {stage084[50]},
      {stage085[48], stage085[49], stage085[50], stage085[51], stage085[52], stage085[53]},
      {stage087[136], stage086[143], stage085[152], stage084[159], stage083[195]}
   );
   gpc1_1 gpc1_1_2798(
      {stage084[51]},
      {stage084[160]}
   );
   gpc1_1 gpc1_1_2799(
      {stage084[52]},
      {stage084[161]}
   );
   gpc1_1 gpc1_1_2800(
      {stage084[53]},
      {stage084[162]}
   );
   gpc1_1 gpc1_1_2801(
      {stage084[54]},
      {stage084[163]}
   );
   gpc1_1 gpc1_1_2802(
      {stage084[55]},
      {stage084[164]}
   );
   gpc1_1 gpc1_1_2803(
      {stage084[56]},
      {stage084[165]}
   );
   gpc1_1 gpc1_1_2804(
      {stage084[57]},
      {stage084[166]}
   );
   gpc1_1 gpc1_1_2805(
      {stage084[58]},
      {stage084[167]}
   );
   gpc1_1 gpc1_1_2806(
      {stage084[59]},
      {stage084[168]}
   );
   gpc1_1 gpc1_1_2807(
      {stage084[60]},
      {stage084[169]}
   );
   gpc1_1 gpc1_1_2808(
      {stage084[61]},
      {stage084[170]}
   );
   gpc1_1 gpc1_1_2809(
      {stage084[62]},
      {stage084[171]}
   );
   gpc1_1 gpc1_1_2810(
      {stage084[63]},
      {stage084[172]}
   );
   gpc1_1 gpc1_1_2811(
      {stage084[64]},
      {stage084[173]}
   );
   gpc1_1 gpc1_1_2812(
      {stage084[65]},
      {stage084[174]}
   );
   gpc1_1 gpc1_1_2813(
      {stage084[66]},
      {stage084[175]}
   );
   gpc1_1 gpc1_1_2814(
      {stage084[67]},
      {stage084[176]}
   );
   gpc1_1 gpc1_1_2815(
      {stage084[68]},
      {stage084[177]}
   );
   gpc1_1 gpc1_1_2816(
      {stage084[69]},
      {stage084[178]}
   );
   gpc1_1 gpc1_1_2817(
      {stage084[70]},
      {stage084[179]}
   );
   gpc1_1 gpc1_1_2818(
      {stage084[71]},
      {stage084[180]}
   );
   gpc1_1 gpc1_1_2819(
      {stage084[72]},
      {stage084[181]}
   );
   gpc1_1 gpc1_1_2820(
      {stage084[73]},
      {stage084[182]}
   );
   gpc1_1 gpc1_1_2821(
      {stage084[74]},
      {stage084[183]}
   );
   gpc1_1 gpc1_1_2822(
      {stage084[75]},
      {stage084[184]}
   );
   gpc1_1 gpc1_1_2823(
      {stage084[76]},
      {stage084[185]}
   );
   gpc1_1 gpc1_1_2824(
      {stage084[77]},
      {stage084[186]}
   );
   gpc606_5 gpc606_5_2825(
      {stage084[78], stage084[79], stage084[80], stage084[81], stage084[82], stage084[83]},
      {stage086[0], stage086[1], stage086[2], stage086[3], stage086[4], stage086[5]},
      {stage088[128], stage087[137], stage086[144], stage085[153], stage084[187]}
   );
   gpc606_5 gpc606_5_2826(
      {stage084[84], stage084[85], stage084[86], stage084[87], stage084[88], stage084[89]},
      {stage086[6], stage086[7], stage086[8], stage086[9], stage086[10], stage086[11]},
      {stage088[129], stage087[138], stage086[145], stage085[154], stage084[188]}
   );
   gpc615_5 gpc615_5_2827(
      {stage084[90], stage084[91], stage084[92], stage084[93], stage084[94]},
      {stage085[54]},
      {stage086[12], stage086[13], stage086[14], stage086[15], stage086[16], stage086[17]},
      {stage088[130], stage087[139], stage086[146], stage085[155], stage084[189]}
   );
   gpc615_5 gpc615_5_2828(
      {stage084[95], stage084[96], stage084[97], stage084[98], stage084[99]},
      {stage085[55]},
      {stage086[18], stage086[19], stage086[20], stage086[21], stage086[22], stage086[23]},
      {stage088[131], stage087[140], stage086[147], stage085[156], stage084[190]}
   );
   gpc615_5 gpc615_5_2829(
      {stage084[100], stage084[101], stage084[102], stage084[103], stage084[104]},
      {stage085[56]},
      {stage086[24], stage086[25], stage086[26], stage086[27], stage086[28], stage086[29]},
      {stage088[132], stage087[141], stage086[148], stage085[157], stage084[191]}
   );
   gpc615_5 gpc615_5_2830(
      {stage084[105], stage084[106], stage084[107], stage084[108], stage084[109]},
      {stage085[57]},
      {stage086[30], stage086[31], stage086[32], stage086[33], stage086[34], stage086[35]},
      {stage088[133], stage087[142], stage086[149], stage085[158], stage084[192]}
   );
   gpc615_5 gpc615_5_2831(
      {stage084[110], stage084[111], stage084[112], stage084[113], stage084[114]},
      {stage085[58]},
      {stage086[36], stage086[37], stage086[38], stage086[39], stage086[40], stage086[41]},
      {stage088[134], stage087[143], stage086[150], stage085[159], stage084[193]}
   );
   gpc615_5 gpc615_5_2832(
      {stage084[115], stage084[116], stage084[117], stage084[118], stage084[119]},
      {stage085[59]},
      {stage086[42], stage086[43], stage086[44], stage086[45], stage086[46], stage086[47]},
      {stage088[135], stage087[144], stage086[151], stage085[160], stage084[194]}
   );
   gpc615_5 gpc615_5_2833(
      {stage084[120], stage084[121], stage084[122], stage084[123], stage084[124]},
      {stage085[60]},
      {stage086[48], stage086[49], stage086[50], stage086[51], stage086[52], stage086[53]},
      {stage088[136], stage087[145], stage086[152], stage085[161], stage084[195]}
   );
   gpc1343_5 gpc1343_5_2834(
      {stage084[125], stage084[126], stage084[127]},
      {stage085[61], stage085[62], stage085[63], stage085[64]},
      {stage086[54], stage086[55], stage086[56]},
      {stage087[0]},
      {stage088[137], stage087[146], stage086[153], stage085[162], stage084[196]}
   );
   gpc1_1 gpc1_1_2835(
      {stage085[65]},
      {stage085[163]}
   );
   gpc1_1 gpc1_1_2836(
      {stage085[66]},
      {stage085[164]}
   );
   gpc1_1 gpc1_1_2837(
      {stage085[67]},
      {stage085[165]}
   );
   gpc1_1 gpc1_1_2838(
      {stage085[68]},
      {stage085[166]}
   );
   gpc1_1 gpc1_1_2839(
      {stage085[69]},
      {stage085[167]}
   );
   gpc1_1 gpc1_1_2840(
      {stage085[70]},
      {stage085[168]}
   );
   gpc1_1 gpc1_1_2841(
      {stage085[71]},
      {stage085[169]}
   );
   gpc1_1 gpc1_1_2842(
      {stage085[72]},
      {stage085[170]}
   );
   gpc1_1 gpc1_1_2843(
      {stage085[73]},
      {stage085[171]}
   );
   gpc1_1 gpc1_1_2844(
      {stage085[74]},
      {stage085[172]}
   );
   gpc1_1 gpc1_1_2845(
      {stage085[75]},
      {stage085[173]}
   );
   gpc1_1 gpc1_1_2846(
      {stage085[76]},
      {stage085[174]}
   );
   gpc1_1 gpc1_1_2847(
      {stage085[77]},
      {stage085[175]}
   );
   gpc1_1 gpc1_1_2848(
      {stage085[78]},
      {stage085[176]}
   );
   gpc1_1 gpc1_1_2849(
      {stage085[79]},
      {stage085[177]}
   );
   gpc1_1 gpc1_1_2850(
      {stage085[80]},
      {stage085[178]}
   );
   gpc1_1 gpc1_1_2851(
      {stage085[81]},
      {stage085[179]}
   );
   gpc1_1 gpc1_1_2852(
      {stage085[82]},
      {stage085[180]}
   );
   gpc1_1 gpc1_1_2853(
      {stage085[83]},
      {stage085[181]}
   );
   gpc1_1 gpc1_1_2854(
      {stage085[84]},
      {stage085[182]}
   );
   gpc1_1 gpc1_1_2855(
      {stage085[85]},
      {stage085[183]}
   );
   gpc1_1 gpc1_1_2856(
      {stage085[86]},
      {stage085[184]}
   );
   gpc1_1 gpc1_1_2857(
      {stage085[87]},
      {stage085[185]}
   );
   gpc1_1 gpc1_1_2858(
      {stage085[88]},
      {stage085[186]}
   );
   gpc1_1 gpc1_1_2859(
      {stage085[89]},
      {stage085[187]}
   );
   gpc1_1 gpc1_1_2860(
      {stage085[90]},
      {stage085[188]}
   );
   gpc1_1 gpc1_1_2861(
      {stage085[91]},
      {stage085[189]}
   );
   gpc1_1 gpc1_1_2862(
      {stage085[92]},
      {stage085[190]}
   );
   gpc1_1 gpc1_1_2863(
      {stage085[93]},
      {stage085[191]}
   );
   gpc1_1 gpc1_1_2864(
      {stage085[94]},
      {stage085[192]}
   );
   gpc1_1 gpc1_1_2865(
      {stage085[95]},
      {stage085[193]}
   );
   gpc1_1 gpc1_1_2866(
      {stage085[96]},
      {stage085[194]}
   );
   gpc1_1 gpc1_1_2867(
      {stage085[97]},
      {stage085[195]}
   );
   gpc1_1 gpc1_1_2868(
      {stage085[98]},
      {stage085[196]}
   );
   gpc1_1 gpc1_1_2869(
      {stage085[99]},
      {stage085[197]}
   );
   gpc1_1 gpc1_1_2870(
      {stage085[100]},
      {stage085[198]}
   );
   gpc1_1 gpc1_1_2871(
      {stage085[101]},
      {stage085[199]}
   );
   gpc1_1 gpc1_1_2872(
      {stage085[102]},
      {stage085[200]}
   );
   gpc1_1 gpc1_1_2873(
      {stage085[103]},
      {stage085[201]}
   );
   gpc1_1 gpc1_1_2874(
      {stage085[104]},
      {stage085[202]}
   );
   gpc1_1 gpc1_1_2875(
      {stage085[105]},
      {stage085[203]}
   );
   gpc1_1 gpc1_1_2876(
      {stage085[106]},
      {stage085[204]}
   );
   gpc1_1 gpc1_1_2877(
      {stage085[107]},
      {stage085[205]}
   );
   gpc1_1 gpc1_1_2878(
      {stage085[108]},
      {stage085[206]}
   );
   gpc1_1 gpc1_1_2879(
      {stage085[109]},
      {stage085[207]}
   );
   gpc1_1 gpc1_1_2880(
      {stage085[110]},
      {stage085[208]}
   );
   gpc1_1 gpc1_1_2881(
      {stage085[111]},
      {stage085[209]}
   );
   gpc1_1 gpc1_1_2882(
      {stage085[112]},
      {stage085[210]}
   );
   gpc1_1 gpc1_1_2883(
      {stage085[113]},
      {stage085[211]}
   );
   gpc1_1 gpc1_1_2884(
      {stage085[114]},
      {stage085[212]}
   );
   gpc1_1 gpc1_1_2885(
      {stage085[115]},
      {stage085[213]}
   );
   gpc1_1 gpc1_1_2886(
      {stage085[116]},
      {stage085[214]}
   );
   gpc1_1 gpc1_1_2887(
      {stage085[117]},
      {stage085[215]}
   );
   gpc615_5 gpc615_5_2888(
      {stage085[118], stage085[119], stage085[120], stage085[121], stage085[122]},
      {stage086[57]},
      {stage087[1], stage087[2], stage087[3], stage087[4], stage087[5], stage087[6]},
      {stage089[128], stage088[138], stage087[147], stage086[154], stage085[216]}
   );
   gpc615_5 gpc615_5_2889(
      {stage085[123], stage085[124], stage085[125], stage085[126], stage085[127]},
      {stage086[58]},
      {stage087[7], stage087[8], stage087[9], stage087[10], stage087[11], stage087[12]},
      {stage089[129], stage088[139], stage087[148], stage086[155], stage085[217]}
   );
   gpc1_1 gpc1_1_2890(
      {stage086[59]},
      {stage086[156]}
   );
   gpc1_1 gpc1_1_2891(
      {stage086[60]},
      {stage086[157]}
   );
   gpc1_1 gpc1_1_2892(
      {stage086[61]},
      {stage086[158]}
   );
   gpc1_1 gpc1_1_2893(
      {stage086[62]},
      {stage086[159]}
   );
   gpc1_1 gpc1_1_2894(
      {stage086[63]},
      {stage086[160]}
   );
   gpc1_1 gpc1_1_2895(
      {stage086[64]},
      {stage086[161]}
   );
   gpc1_1 gpc1_1_2896(
      {stage086[65]},
      {stage086[162]}
   );
   gpc1_1 gpc1_1_2897(
      {stage086[66]},
      {stage086[163]}
   );
   gpc1_1 gpc1_1_2898(
      {stage086[67]},
      {stage086[164]}
   );
   gpc1_1 gpc1_1_2899(
      {stage086[68]},
      {stage086[165]}
   );
   gpc1_1 gpc1_1_2900(
      {stage086[69]},
      {stage086[166]}
   );
   gpc1_1 gpc1_1_2901(
      {stage086[70]},
      {stage086[167]}
   );
   gpc1_1 gpc1_1_2902(
      {stage086[71]},
      {stage086[168]}
   );
   gpc1_1 gpc1_1_2903(
      {stage086[72]},
      {stage086[169]}
   );
   gpc1_1 gpc1_1_2904(
      {stage086[73]},
      {stage086[170]}
   );
   gpc1_1 gpc1_1_2905(
      {stage086[74]},
      {stage086[171]}
   );
   gpc1_1 gpc1_1_2906(
      {stage086[75]},
      {stage086[172]}
   );
   gpc1_1 gpc1_1_2907(
      {stage086[76]},
      {stage086[173]}
   );
   gpc1_1 gpc1_1_2908(
      {stage086[77]},
      {stage086[174]}
   );
   gpc1_1 gpc1_1_2909(
      {stage086[78]},
      {stage086[175]}
   );
   gpc1_1 gpc1_1_2910(
      {stage086[79]},
      {stage086[176]}
   );
   gpc1_1 gpc1_1_2911(
      {stage086[80]},
      {stage086[177]}
   );
   gpc1_1 gpc1_1_2912(
      {stage086[81]},
      {stage086[178]}
   );
   gpc1_1 gpc1_1_2913(
      {stage086[82]},
      {stage086[179]}
   );
   gpc1_1 gpc1_1_2914(
      {stage086[83]},
      {stage086[180]}
   );
   gpc1_1 gpc1_1_2915(
      {stage086[84]},
      {stage086[181]}
   );
   gpc1_1 gpc1_1_2916(
      {stage086[85]},
      {stage086[182]}
   );
   gpc1_1 gpc1_1_2917(
      {stage086[86]},
      {stage086[183]}
   );
   gpc1_1 gpc1_1_2918(
      {stage086[87]},
      {stage086[184]}
   );
   gpc1_1 gpc1_1_2919(
      {stage086[88]},
      {stage086[185]}
   );
   gpc1_1 gpc1_1_2920(
      {stage086[89]},
      {stage086[186]}
   );
   gpc1_1 gpc1_1_2921(
      {stage086[90]},
      {stage086[187]}
   );
   gpc1_1 gpc1_1_2922(
      {stage086[91]},
      {stage086[188]}
   );
   gpc1_1 gpc1_1_2923(
      {stage086[92]},
      {stage086[189]}
   );
   gpc1_1 gpc1_1_2924(
      {stage086[93]},
      {stage086[190]}
   );
   gpc1_1 gpc1_1_2925(
      {stage086[94]},
      {stage086[191]}
   );
   gpc1_1 gpc1_1_2926(
      {stage086[95]},
      {stage086[192]}
   );
   gpc1_1 gpc1_1_2927(
      {stage086[96]},
      {stage086[193]}
   );
   gpc1_1 gpc1_1_2928(
      {stage086[97]},
      {stage086[194]}
   );
   gpc1_1 gpc1_1_2929(
      {stage086[98]},
      {stage086[195]}
   );
   gpc1_1 gpc1_1_2930(
      {stage086[99]},
      {stage086[196]}
   );
   gpc1_1 gpc1_1_2931(
      {stage086[100]},
      {stage086[197]}
   );
   gpc1_1 gpc1_1_2932(
      {stage086[101]},
      {stage086[198]}
   );
   gpc1_1 gpc1_1_2933(
      {stage086[102]},
      {stage086[199]}
   );
   gpc1_1 gpc1_1_2934(
      {stage086[103]},
      {stage086[200]}
   );
   gpc606_5 gpc606_5_2935(
      {stage086[104], stage086[105], stage086[106], stage086[107], stage086[108], stage086[109]},
      {stage088[0], stage088[1], stage088[2], stage088[3], stage088[4], stage088[5]},
      {stage090[128], stage089[130], stage088[140], stage087[149], stage086[201]}
   );
   gpc606_5 gpc606_5_2936(
      {stage086[110], stage086[111], stage086[112], stage086[113], stage086[114], stage086[115]},
      {stage088[6], stage088[7], stage088[8], stage088[9], stage088[10], stage088[11]},
      {stage090[129], stage089[131], stage088[141], stage087[150], stage086[202]}
   );
   gpc606_5 gpc606_5_2937(
      {stage086[116], stage086[117], stage086[118], stage086[119], stage086[120], stage086[121]},
      {stage088[12], stage088[13], stage088[14], stage088[15], stage088[16], stage088[17]},
      {stage090[130], stage089[132], stage088[142], stage087[151], stage086[203]}
   );
   gpc606_5 gpc606_5_2938(
      {stage086[122], stage086[123], stage086[124], stage086[125], stage086[126], stage086[127]},
      {stage088[18], stage088[19], stage088[20], stage088[21], stage088[22], stage088[23]},
      {stage090[131], stage089[133], stage088[143], stage087[152], stage086[204]}
   );
   gpc1_1 gpc1_1_2939(
      {stage087[13]},
      {stage087[153]}
   );
   gpc1_1 gpc1_1_2940(
      {stage087[14]},
      {stage087[154]}
   );
   gpc1_1 gpc1_1_2941(
      {stage087[15]},
      {stage087[155]}
   );
   gpc1_1 gpc1_1_2942(
      {stage087[16]},
      {stage087[156]}
   );
   gpc1_1 gpc1_1_2943(
      {stage087[17]},
      {stage087[157]}
   );
   gpc1_1 gpc1_1_2944(
      {stage087[18]},
      {stage087[158]}
   );
   gpc1_1 gpc1_1_2945(
      {stage087[19]},
      {stage087[159]}
   );
   gpc1_1 gpc1_1_2946(
      {stage087[20]},
      {stage087[160]}
   );
   gpc1_1 gpc1_1_2947(
      {stage087[21]},
      {stage087[161]}
   );
   gpc1_1 gpc1_1_2948(
      {stage087[22]},
      {stage087[162]}
   );
   gpc1_1 gpc1_1_2949(
      {stage087[23]},
      {stage087[163]}
   );
   gpc1_1 gpc1_1_2950(
      {stage087[24]},
      {stage087[164]}
   );
   gpc1_1 gpc1_1_2951(
      {stage087[25]},
      {stage087[165]}
   );
   gpc606_5 gpc606_5_2952(
      {stage087[26], stage087[27], stage087[28], stage087[29], stage087[30], stage087[31]},
      {stage089[0], stage089[1], stage089[2], stage089[3], stage089[4], stage089[5]},
      {stage091[128], stage090[132], stage089[134], stage088[144], stage087[166]}
   );
   gpc606_5 gpc606_5_2953(
      {stage087[32], stage087[33], stage087[34], stage087[35], stage087[36], stage087[37]},
      {stage089[6], stage089[7], stage089[8], stage089[9], stage089[10], stage089[11]},
      {stage091[129], stage090[133], stage089[135], stage088[145], stage087[167]}
   );
   gpc606_5 gpc606_5_2954(
      {stage087[38], stage087[39], stage087[40], stage087[41], stage087[42], stage087[43]},
      {stage089[12], stage089[13], stage089[14], stage089[15], stage089[16], stage089[17]},
      {stage091[130], stage090[134], stage089[136], stage088[146], stage087[168]}
   );
   gpc606_5 gpc606_5_2955(
      {stage087[44], stage087[45], stage087[46], stage087[47], stage087[48], stage087[49]},
      {stage089[18], stage089[19], stage089[20], stage089[21], stage089[22], stage089[23]},
      {stage091[131], stage090[135], stage089[137], stage088[147], stage087[169]}
   );
   gpc606_5 gpc606_5_2956(
      {stage087[50], stage087[51], stage087[52], stage087[53], stage087[54], stage087[55]},
      {stage089[24], stage089[25], stage089[26], stage089[27], stage089[28], stage089[29]},
      {stage091[132], stage090[136], stage089[138], stage088[148], stage087[170]}
   );
   gpc606_5 gpc606_5_2957(
      {stage087[56], stage087[57], stage087[58], stage087[59], stage087[60], stage087[61]},
      {stage089[30], stage089[31], stage089[32], stage089[33], stage089[34], stage089[35]},
      {stage091[133], stage090[137], stage089[139], stage088[149], stage087[171]}
   );
   gpc606_5 gpc606_5_2958(
      {stage087[62], stage087[63], stage087[64], stage087[65], stage087[66], stage087[67]},
      {stage089[36], stage089[37], stage089[38], stage089[39], stage089[40], stage089[41]},
      {stage091[134], stage090[138], stage089[140], stage088[150], stage087[172]}
   );
   gpc606_5 gpc606_5_2959(
      {stage087[68], stage087[69], stage087[70], stage087[71], stage087[72], stage087[73]},
      {stage089[42], stage089[43], stage089[44], stage089[45], stage089[46], stage089[47]},
      {stage091[135], stage090[139], stage089[141], stage088[151], stage087[173]}
   );
   gpc606_5 gpc606_5_2960(
      {stage087[74], stage087[75], stage087[76], stage087[77], stage087[78], stage087[79]},
      {stage089[48], stage089[49], stage089[50], stage089[51], stage089[52], stage089[53]},
      {stage091[136], stage090[140], stage089[142], stage088[152], stage087[174]}
   );
   gpc606_5 gpc606_5_2961(
      {stage087[80], stage087[81], stage087[82], stage087[83], stage087[84], stage087[85]},
      {stage089[54], stage089[55], stage089[56], stage089[57], stage089[58], stage089[59]},
      {stage091[137], stage090[141], stage089[143], stage088[153], stage087[175]}
   );
   gpc606_5 gpc606_5_2962(
      {stage087[86], stage087[87], stage087[88], stage087[89], stage087[90], stage087[91]},
      {stage089[60], stage089[61], stage089[62], stage089[63], stage089[64], stage089[65]},
      {stage091[138], stage090[142], stage089[144], stage088[154], stage087[176]}
   );
   gpc606_5 gpc606_5_2963(
      {stage087[92], stage087[93], stage087[94], stage087[95], stage087[96], stage087[97]},
      {stage089[66], stage089[67], stage089[68], stage089[69], stage089[70], stage089[71]},
      {stage091[139], stage090[143], stage089[145], stage088[155], stage087[177]}
   );
   gpc606_5 gpc606_5_2964(
      {stage087[98], stage087[99], stage087[100], stage087[101], stage087[102], stage087[103]},
      {stage089[72], stage089[73], stage089[74], stage089[75], stage089[76], stage089[77]},
      {stage091[140], stage090[144], stage089[146], stage088[156], stage087[178]}
   );
   gpc606_5 gpc606_5_2965(
      {stage087[104], stage087[105], stage087[106], stage087[107], stage087[108], stage087[109]},
      {stage089[78], stage089[79], stage089[80], stage089[81], stage089[82], stage089[83]},
      {stage091[141], stage090[145], stage089[147], stage088[157], stage087[179]}
   );
   gpc606_5 gpc606_5_2966(
      {stage087[110], stage087[111], stage087[112], stage087[113], stage087[114], stage087[115]},
      {stage089[84], stage089[85], stage089[86], stage089[87], stage089[88], stage089[89]},
      {stage091[142], stage090[146], stage089[148], stage088[158], stage087[180]}
   );
   gpc606_5 gpc606_5_2967(
      {stage087[116], stage087[117], stage087[118], stage087[119], stage087[120], stage087[121]},
      {stage089[90], stage089[91], stage089[92], stage089[93], stage089[94], stage089[95]},
      {stage091[143], stage090[147], stage089[149], stage088[159], stage087[181]}
   );
   gpc606_5 gpc606_5_2968(
      {stage087[122], stage087[123], stage087[124], stage087[125], stage087[126], stage087[127]},
      {stage089[96], stage089[97], stage089[98], stage089[99], stage089[100], stage089[101]},
      {stage091[144], stage090[148], stage089[150], stage088[160], stage087[182]}
   );
   gpc1_1 gpc1_1_2969(
      {stage088[24]},
      {stage088[161]}
   );
   gpc1_1 gpc1_1_2970(
      {stage088[25]},
      {stage088[162]}
   );
   gpc1_1 gpc1_1_2971(
      {stage088[26]},
      {stage088[163]}
   );
   gpc1_1 gpc1_1_2972(
      {stage088[27]},
      {stage088[164]}
   );
   gpc1_1 gpc1_1_2973(
      {stage088[28]},
      {stage088[165]}
   );
   gpc1_1 gpc1_1_2974(
      {stage088[29]},
      {stage088[166]}
   );
   gpc1_1 gpc1_1_2975(
      {stage088[30]},
      {stage088[167]}
   );
   gpc1_1 gpc1_1_2976(
      {stage088[31]},
      {stage088[168]}
   );
   gpc1_1 gpc1_1_2977(
      {stage088[32]},
      {stage088[169]}
   );
   gpc1_1 gpc1_1_2978(
      {stage088[33]},
      {stage088[170]}
   );
   gpc1_1 gpc1_1_2979(
      {stage088[34]},
      {stage088[171]}
   );
   gpc1_1 gpc1_1_2980(
      {stage088[35]},
      {stage088[172]}
   );
   gpc1_1 gpc1_1_2981(
      {stage088[36]},
      {stage088[173]}
   );
   gpc1_1 gpc1_1_2982(
      {stage088[37]},
      {stage088[174]}
   );
   gpc1_1 gpc1_1_2983(
      {stage088[38]},
      {stage088[175]}
   );
   gpc1_1 gpc1_1_2984(
      {stage088[39]},
      {stage088[176]}
   );
   gpc1_1 gpc1_1_2985(
      {stage088[40]},
      {stage088[177]}
   );
   gpc1_1 gpc1_1_2986(
      {stage088[41]},
      {stage088[178]}
   );
   gpc1_1 gpc1_1_2987(
      {stage088[42]},
      {stage088[179]}
   );
   gpc1_1 gpc1_1_2988(
      {stage088[43]},
      {stage088[180]}
   );
   gpc1_1 gpc1_1_2989(
      {stage088[44]},
      {stage088[181]}
   );
   gpc1_1 gpc1_1_2990(
      {stage088[45]},
      {stage088[182]}
   );
   gpc1_1 gpc1_1_2991(
      {stage088[46]},
      {stage088[183]}
   );
   gpc1_1 gpc1_1_2992(
      {stage088[47]},
      {stage088[184]}
   );
   gpc1_1 gpc1_1_2993(
      {stage088[48]},
      {stage088[185]}
   );
   gpc1_1 gpc1_1_2994(
      {stage088[49]},
      {stage088[186]}
   );
   gpc1_1 gpc1_1_2995(
      {stage088[50]},
      {stage088[187]}
   );
   gpc1_1 gpc1_1_2996(
      {stage088[51]},
      {stage088[188]}
   );
   gpc1_1 gpc1_1_2997(
      {stage088[52]},
      {stage088[189]}
   );
   gpc1_1 gpc1_1_2998(
      {stage088[53]},
      {stage088[190]}
   );
   gpc1_1 gpc1_1_2999(
      {stage088[54]},
      {stage088[191]}
   );
   gpc1_1 gpc1_1_3000(
      {stage088[55]},
      {stage088[192]}
   );
   gpc1_1 gpc1_1_3001(
      {stage088[56]},
      {stage088[193]}
   );
   gpc1_1 gpc1_1_3002(
      {stage088[57]},
      {stage088[194]}
   );
   gpc1_1 gpc1_1_3003(
      {stage088[58]},
      {stage088[195]}
   );
   gpc1_1 gpc1_1_3004(
      {stage088[59]},
      {stage088[196]}
   );
   gpc1_1 gpc1_1_3005(
      {stage088[60]},
      {stage088[197]}
   );
   gpc1_1 gpc1_1_3006(
      {stage088[61]},
      {stage088[198]}
   );
   gpc1_1 gpc1_1_3007(
      {stage088[62]},
      {stage088[199]}
   );
   gpc1_1 gpc1_1_3008(
      {stage088[63]},
      {stage088[200]}
   );
   gpc1_1 gpc1_1_3009(
      {stage088[64]},
      {stage088[201]}
   );
   gpc1_1 gpc1_1_3010(
      {stage088[65]},
      {stage088[202]}
   );
   gpc1_1 gpc1_1_3011(
      {stage088[66]},
      {stage088[203]}
   );
   gpc1_1 gpc1_1_3012(
      {stage088[67]},
      {stage088[204]}
   );
   gpc1_1 gpc1_1_3013(
      {stage088[68]},
      {stage088[205]}
   );
   gpc1_1 gpc1_1_3014(
      {stage088[69]},
      {stage088[206]}
   );
   gpc1_1 gpc1_1_3015(
      {stage088[70]},
      {stage088[207]}
   );
   gpc1_1 gpc1_1_3016(
      {stage088[71]},
      {stage088[208]}
   );
   gpc1_1 gpc1_1_3017(
      {stage088[72]},
      {stage088[209]}
   );
   gpc1_1 gpc1_1_3018(
      {stage088[73]},
      {stage088[210]}
   );
   gpc606_5 gpc606_5_3019(
      {stage088[74], stage088[75], stage088[76], stage088[77], stage088[78], stage088[79]},
      {stage090[0], stage090[1], stage090[2], stage090[3], stage090[4], stage090[5]},
      {stage092[128], stage091[145], stage090[149], stage089[151], stage088[211]}
   );
   gpc606_5 gpc606_5_3020(
      {stage088[80], stage088[81], stage088[82], stage088[83], stage088[84], stage088[85]},
      {stage090[6], stage090[7], stage090[8], stage090[9], stage090[10], stage090[11]},
      {stage092[129], stage091[146], stage090[150], stage089[152], stage088[212]}
   );
   gpc606_5 gpc606_5_3021(
      {stage088[86], stage088[87], stage088[88], stage088[89], stage088[90], stage088[91]},
      {stage090[12], stage090[13], stage090[14], stage090[15], stage090[16], stage090[17]},
      {stage092[130], stage091[147], stage090[151], stage089[153], stage088[213]}
   );
   gpc606_5 gpc606_5_3022(
      {stage088[92], stage088[93], stage088[94], stage088[95], stage088[96], stage088[97]},
      {stage090[18], stage090[19], stage090[20], stage090[21], stage090[22], stage090[23]},
      {stage092[131], stage091[148], stage090[152], stage089[154], stage088[214]}
   );
   gpc606_5 gpc606_5_3023(
      {stage088[98], stage088[99], stage088[100], stage088[101], stage088[102], stage088[103]},
      {stage090[24], stage090[25], stage090[26], stage090[27], stage090[28], stage090[29]},
      {stage092[132], stage091[149], stage090[153], stage089[155], stage088[215]}
   );
   gpc606_5 gpc606_5_3024(
      {stage088[104], stage088[105], stage088[106], stage088[107], stage088[108], stage088[109]},
      {stage090[30], stage090[31], stage090[32], stage090[33], stage090[34], stage090[35]},
      {stage092[133], stage091[150], stage090[154], stage089[156], stage088[216]}
   );
   gpc606_5 gpc606_5_3025(
      {stage088[110], stage088[111], stage088[112], stage088[113], stage088[114], stage088[115]},
      {stage090[36], stage090[37], stage090[38], stage090[39], stage090[40], stage090[41]},
      {stage092[134], stage091[151], stage090[155], stage089[157], stage088[217]}
   );
   gpc606_5 gpc606_5_3026(
      {stage088[116], stage088[117], stage088[118], stage088[119], stage088[120], stage088[121]},
      {stage090[42], stage090[43], stage090[44], stage090[45], stage090[46], stage090[47]},
      {stage092[135], stage091[152], stage090[156], stage089[158], stage088[218]}
   );
   gpc606_5 gpc606_5_3027(
      {stage088[122], stage088[123], stage088[124], stage088[125], stage088[126], stage088[127]},
      {stage090[48], stage090[49], stage090[50], stage090[51], stage090[52], stage090[53]},
      {stage092[136], stage091[153], stage090[157], stage089[159], stage088[219]}
   );
   gpc1_1 gpc1_1_3028(
      {stage089[102]},
      {stage089[160]}
   );
   gpc615_5 gpc615_5_3029(
      {stage089[103], stage089[104], stage089[105], stage089[106], stage089[107]},
      {stage090[54]},
      {stage091[0], stage091[1], stage091[2], stage091[3], stage091[4], stage091[5]},
      {stage093[128], stage092[137], stage091[154], stage090[158], stage089[161]}
   );
   gpc615_5 gpc615_5_3030(
      {stage089[108], stage089[109], stage089[110], stage089[111], stage089[112]},
      {stage090[55]},
      {stage091[6], stage091[7], stage091[8], stage091[9], stage091[10], stage091[11]},
      {stage093[129], stage092[138], stage091[155], stage090[159], stage089[162]}
   );
   gpc615_5 gpc615_5_3031(
      {stage089[113], stage089[114], stage089[115], stage089[116], stage089[117]},
      {stage090[56]},
      {stage091[12], stage091[13], stage091[14], stage091[15], stage091[16], stage091[17]},
      {stage093[130], stage092[139], stage091[156], stage090[160], stage089[163]}
   );
   gpc615_5 gpc615_5_3032(
      {stage089[118], stage089[119], stage089[120], stage089[121], stage089[122]},
      {stage090[57]},
      {stage091[18], stage091[19], stage091[20], stage091[21], stage091[22], stage091[23]},
      {stage093[131], stage092[140], stage091[157], stage090[161], stage089[164]}
   );
   gpc615_5 gpc615_5_3033(
      {stage089[123], stage089[124], stage089[125], stage089[126], stage089[127]},
      {stage090[58]},
      {stage091[24], stage091[25], stage091[26], stage091[27], stage091[28], stage091[29]},
      {stage093[132], stage092[141], stage091[158], stage090[162], stage089[165]}
   );
   gpc1_1 gpc1_1_3034(
      {stage090[59]},
      {stage090[163]}
   );
   gpc1_1 gpc1_1_3035(
      {stage090[60]},
      {stage090[164]}
   );
   gpc1_1 gpc1_1_3036(
      {stage090[61]},
      {stage090[165]}
   );
   gpc1_1 gpc1_1_3037(
      {stage090[62]},
      {stage090[166]}
   );
   gpc1_1 gpc1_1_3038(
      {stage090[63]},
      {stage090[167]}
   );
   gpc1_1 gpc1_1_3039(
      {stage090[64]},
      {stage090[168]}
   );
   gpc606_5 gpc606_5_3040(
      {stage090[65], stage090[66], stage090[67], stage090[68], stage090[69], stage090[70]},
      {stage092[0], stage092[1], stage092[2], stage092[3], stage092[4], stage092[5]},
      {stage094[128], stage093[133], stage092[142], stage091[159], stage090[169]}
   );
   gpc606_5 gpc606_5_3041(
      {stage090[71], stage090[72], stage090[73], stage090[74], stage090[75], stage090[76]},
      {stage092[6], stage092[7], stage092[8], stage092[9], stage092[10], stage092[11]},
      {stage094[129], stage093[134], stage092[143], stage091[160], stage090[170]}
   );
   gpc606_5 gpc606_5_3042(
      {stage090[77], stage090[78], stage090[79], stage090[80], stage090[81], stage090[82]},
      {stage092[12], stage092[13], stage092[14], stage092[15], stage092[16], stage092[17]},
      {stage094[130], stage093[135], stage092[144], stage091[161], stage090[171]}
   );
   gpc606_5 gpc606_5_3043(
      {stage090[83], stage090[84], stage090[85], stage090[86], stage090[87], stage090[88]},
      {stage092[18], stage092[19], stage092[20], stage092[21], stage092[22], stage092[23]},
      {stage094[131], stage093[136], stage092[145], stage091[162], stage090[172]}
   );
   gpc606_5 gpc606_5_3044(
      {stage090[89], stage090[90], stage090[91], stage090[92], stage090[93], stage090[94]},
      {stage092[24], stage092[25], stage092[26], stage092[27], stage092[28], stage092[29]},
      {stage094[132], stage093[137], stage092[146], stage091[163], stage090[173]}
   );
   gpc606_5 gpc606_5_3045(
      {stage090[95], stage090[96], stage090[97], stage090[98], stage090[99], stage090[100]},
      {stage092[30], stage092[31], stage092[32], stage092[33], stage092[34], stage092[35]},
      {stage094[133], stage093[138], stage092[147], stage091[164], stage090[174]}
   );
   gpc606_5 gpc606_5_3046(
      {stage090[101], stage090[102], stage090[103], stage090[104], stage090[105], stage090[106]},
      {stage092[36], stage092[37], stage092[38], stage092[39], stage092[40], stage092[41]},
      {stage094[134], stage093[139], stage092[148], stage091[165], stage090[175]}
   );
   gpc606_5 gpc606_5_3047(
      {stage090[107], stage090[108], stage090[109], stage090[110], stage090[111], stage090[112]},
      {stage092[42], stage092[43], stage092[44], stage092[45], stage092[46], stage092[47]},
      {stage094[135], stage093[140], stage092[149], stage091[166], stage090[176]}
   );
   gpc615_5 gpc615_5_3048(
      {stage090[113], stage090[114], stage090[115], stage090[116], stage090[117]},
      {stage091[30]},
      {stage092[48], stage092[49], stage092[50], stage092[51], stage092[52], stage092[53]},
      {stage094[136], stage093[141], stage092[150], stage091[167], stage090[177]}
   );
   gpc615_5 gpc615_5_3049(
      {stage090[118], stage090[119], stage090[120], stage090[121], stage090[122]},
      {stage091[31]},
      {stage092[54], stage092[55], stage092[56], stage092[57], stage092[58], stage092[59]},
      {stage094[137], stage093[142], stage092[151], stage091[168], stage090[178]}
   );
   gpc615_5 gpc615_5_3050(
      {stage090[123], stage090[124], stage090[125], stage090[126], stage090[127]},
      {stage091[32]},
      {stage092[60], stage092[61], stage092[62], stage092[63], stage092[64], stage092[65]},
      {stage094[138], stage093[143], stage092[152], stage091[169], stage090[179]}
   );
   gpc1_1 gpc1_1_3051(
      {stage091[33]},
      {stage091[170]}
   );
   gpc1_1 gpc1_1_3052(
      {stage091[34]},
      {stage091[171]}
   );
   gpc1_1 gpc1_1_3053(
      {stage091[35]},
      {stage091[172]}
   );
   gpc1_1 gpc1_1_3054(
      {stage091[36]},
      {stage091[173]}
   );
   gpc1_1 gpc1_1_3055(
      {stage091[37]},
      {stage091[174]}
   );
   gpc1_1 gpc1_1_3056(
      {stage091[38]},
      {stage091[175]}
   );
   gpc1_1 gpc1_1_3057(
      {stage091[39]},
      {stage091[176]}
   );
   gpc1_1 gpc1_1_3058(
      {stage091[40]},
      {stage091[177]}
   );
   gpc1_1 gpc1_1_3059(
      {stage091[41]},
      {stage091[178]}
   );
   gpc1_1 gpc1_1_3060(
      {stage091[42]},
      {stage091[179]}
   );
   gpc1_1 gpc1_1_3061(
      {stage091[43]},
      {stage091[180]}
   );
   gpc1_1 gpc1_1_3062(
      {stage091[44]},
      {stage091[181]}
   );
   gpc1_1 gpc1_1_3063(
      {stage091[45]},
      {stage091[182]}
   );
   gpc1_1 gpc1_1_3064(
      {stage091[46]},
      {stage091[183]}
   );
   gpc1_1 gpc1_1_3065(
      {stage091[47]},
      {stage091[184]}
   );
   gpc1_1 gpc1_1_3066(
      {stage091[48]},
      {stage091[185]}
   );
   gpc1_1 gpc1_1_3067(
      {stage091[49]},
      {stage091[186]}
   );
   gpc606_5 gpc606_5_3068(
      {stage091[50], stage091[51], stage091[52], stage091[53], stage091[54], stage091[55]},
      {stage093[0], stage093[1], stage093[2], stage093[3], stage093[4], stage093[5]},
      {stage095[128], stage094[139], stage093[144], stage092[153], stage091[187]}
   );
   gpc606_5 gpc606_5_3069(
      {stage091[56], stage091[57], stage091[58], stage091[59], stage091[60], stage091[61]},
      {stage093[6], stage093[7], stage093[8], stage093[9], stage093[10], stage093[11]},
      {stage095[129], stage094[140], stage093[145], stage092[154], stage091[188]}
   );
   gpc606_5 gpc606_5_3070(
      {stage091[62], stage091[63], stage091[64], stage091[65], stage091[66], stage091[67]},
      {stage093[12], stage093[13], stage093[14], stage093[15], stage093[16], stage093[17]},
      {stage095[130], stage094[141], stage093[146], stage092[155], stage091[189]}
   );
   gpc606_5 gpc606_5_3071(
      {stage091[68], stage091[69], stage091[70], stage091[71], stage091[72], stage091[73]},
      {stage093[18], stage093[19], stage093[20], stage093[21], stage093[22], stage093[23]},
      {stage095[131], stage094[142], stage093[147], stage092[156], stage091[190]}
   );
   gpc606_5 gpc606_5_3072(
      {stage091[74], stage091[75], stage091[76], stage091[77], stage091[78], stage091[79]},
      {stage093[24], stage093[25], stage093[26], stage093[27], stage093[28], stage093[29]},
      {stage095[132], stage094[143], stage093[148], stage092[157], stage091[191]}
   );
   gpc606_5 gpc606_5_3073(
      {stage091[80], stage091[81], stage091[82], stage091[83], stage091[84], stage091[85]},
      {stage093[30], stage093[31], stage093[32], stage093[33], stage093[34], stage093[35]},
      {stage095[133], stage094[144], stage093[149], stage092[158], stage091[192]}
   );
   gpc606_5 gpc606_5_3074(
      {stage091[86], stage091[87], stage091[88], stage091[89], stage091[90], stage091[91]},
      {stage093[36], stage093[37], stage093[38], stage093[39], stage093[40], stage093[41]},
      {stage095[134], stage094[145], stage093[150], stage092[159], stage091[193]}
   );
   gpc606_5 gpc606_5_3075(
      {stage091[92], stage091[93], stage091[94], stage091[95], stage091[96], stage091[97]},
      {stage093[42], stage093[43], stage093[44], stage093[45], stage093[46], stage093[47]},
      {stage095[135], stage094[146], stage093[151], stage092[160], stage091[194]}
   );
   gpc606_5 gpc606_5_3076(
      {stage091[98], stage091[99], stage091[100], stage091[101], stage091[102], stage091[103]},
      {stage093[48], stage093[49], stage093[50], stage093[51], stage093[52], stage093[53]},
      {stage095[136], stage094[147], stage093[152], stage092[161], stage091[195]}
   );
   gpc606_5 gpc606_5_3077(
      {stage091[104], stage091[105], stage091[106], stage091[107], stage091[108], stage091[109]},
      {stage093[54], stage093[55], stage093[56], stage093[57], stage093[58], stage093[59]},
      {stage095[137], stage094[148], stage093[153], stage092[162], stage091[196]}
   );
   gpc606_5 gpc606_5_3078(
      {stage091[110], stage091[111], stage091[112], stage091[113], stage091[114], stage091[115]},
      {stage093[60], stage093[61], stage093[62], stage093[63], stage093[64], stage093[65]},
      {stage095[138], stage094[149], stage093[154], stage092[163], stage091[197]}
   );
   gpc606_5 gpc606_5_3079(
      {stage091[116], stage091[117], stage091[118], stage091[119], stage091[120], stage091[121]},
      {stage093[66], stage093[67], stage093[68], stage093[69], stage093[70], stage093[71]},
      {stage095[139], stage094[150], stage093[155], stage092[164], stage091[198]}
   );
   gpc606_5 gpc606_5_3080(
      {stage091[122], stage091[123], stage091[124], stage091[125], stage091[126], stage091[127]},
      {stage093[72], stage093[73], stage093[74], stage093[75], stage093[76], stage093[77]},
      {stage095[140], stage094[151], stage093[156], stage092[165], stage091[199]}
   );
   gpc1_1 gpc1_1_3081(
      {stage092[66]},
      {stage092[166]}
   );
   gpc1_1 gpc1_1_3082(
      {stage092[67]},
      {stage092[167]}
   );
   gpc1_1 gpc1_1_3083(
      {stage092[68]},
      {stage092[168]}
   );
   gpc1_1 gpc1_1_3084(
      {stage092[69]},
      {stage092[169]}
   );
   gpc1_1 gpc1_1_3085(
      {stage092[70]},
      {stage092[170]}
   );
   gpc1_1 gpc1_1_3086(
      {stage092[71]},
      {stage092[171]}
   );
   gpc1_1 gpc1_1_3087(
      {stage092[72]},
      {stage092[172]}
   );
   gpc1_1 gpc1_1_3088(
      {stage092[73]},
      {stage092[173]}
   );
   gpc1_1 gpc1_1_3089(
      {stage092[74]},
      {stage092[174]}
   );
   gpc1_1 gpc1_1_3090(
      {stage092[75]},
      {stage092[175]}
   );
   gpc1_1 gpc1_1_3091(
      {stage092[76]},
      {stage092[176]}
   );
   gpc1_1 gpc1_1_3092(
      {stage092[77]},
      {stage092[177]}
   );
   gpc1_1 gpc1_1_3093(
      {stage092[78]},
      {stage092[178]}
   );
   gpc1_1 gpc1_1_3094(
      {stage092[79]},
      {stage092[179]}
   );
   gpc1_1 gpc1_1_3095(
      {stage092[80]},
      {stage092[180]}
   );
   gpc1_1 gpc1_1_3096(
      {stage092[81]},
      {stage092[181]}
   );
   gpc1_1 gpc1_1_3097(
      {stage092[82]},
      {stage092[182]}
   );
   gpc1_1 gpc1_1_3098(
      {stage092[83]},
      {stage092[183]}
   );
   gpc1_1 gpc1_1_3099(
      {stage092[84]},
      {stage092[184]}
   );
   gpc1_1 gpc1_1_3100(
      {stage092[85]},
      {stage092[185]}
   );
   gpc1_1 gpc1_1_3101(
      {stage092[86]},
      {stage092[186]}
   );
   gpc1_1 gpc1_1_3102(
      {stage092[87]},
      {stage092[187]}
   );
   gpc1_1 gpc1_1_3103(
      {stage092[88]},
      {stage092[188]}
   );
   gpc1_1 gpc1_1_3104(
      {stage092[89]},
      {stage092[189]}
   );
   gpc1_1 gpc1_1_3105(
      {stage092[90]},
      {stage092[190]}
   );
   gpc606_5 gpc606_5_3106(
      {stage092[91], stage092[92], stage092[93], stage092[94], stage092[95], stage092[96]},
      {stage094[0], stage094[1], stage094[2], stage094[3], stage094[4], stage094[5]},
      {stage096[128], stage095[141], stage094[152], stage093[157], stage092[191]}
   );
   gpc606_5 gpc606_5_3107(
      {stage092[97], stage092[98], stage092[99], stage092[100], stage092[101], stage092[102]},
      {stage094[6], stage094[7], stage094[8], stage094[9], stage094[10], stage094[11]},
      {stage096[129], stage095[142], stage094[153], stage093[158], stage092[192]}
   );
   gpc615_5 gpc615_5_3108(
      {stage092[103], stage092[104], stage092[105], stage092[106], stage092[107]},
      {stage093[78]},
      {stage094[12], stage094[13], stage094[14], stage094[15], stage094[16], stage094[17]},
      {stage096[130], stage095[143], stage094[154], stage093[159], stage092[193]}
   );
   gpc615_5 gpc615_5_3109(
      {stage092[108], stage092[109], stage092[110], stage092[111], stage092[112]},
      {stage093[79]},
      {stage094[18], stage094[19], stage094[20], stage094[21], stage094[22], stage094[23]},
      {stage096[131], stage095[144], stage094[155], stage093[160], stage092[194]}
   );
   gpc615_5 gpc615_5_3110(
      {stage092[113], stage092[114], stage092[115], stage092[116], stage092[117]},
      {stage093[80]},
      {stage094[24], stage094[25], stage094[26], stage094[27], stage094[28], stage094[29]},
      {stage096[132], stage095[145], stage094[156], stage093[161], stage092[195]}
   );
   gpc615_5 gpc615_5_3111(
      {stage092[118], stage092[119], stage092[120], stage092[121], stage092[122]},
      {stage093[81]},
      {stage094[30], stage094[31], stage094[32], stage094[33], stage094[34], stage094[35]},
      {stage096[133], stage095[146], stage094[157], stage093[162], stage092[196]}
   );
   gpc615_5 gpc615_5_3112(
      {stage092[123], stage092[124], stage092[125], stage092[126], stage092[127]},
      {stage093[82]},
      {stage094[36], stage094[37], stage094[38], stage094[39], stage094[40], stage094[41]},
      {stage096[134], stage095[147], stage094[158], stage093[163], stage092[197]}
   );
   gpc1_1 gpc1_1_3113(
      {stage093[83]},
      {stage093[164]}
   );
   gpc1_1 gpc1_1_3114(
      {stage093[84]},
      {stage093[165]}
   );
   gpc1_1 gpc1_1_3115(
      {stage093[85]},
      {stage093[166]}
   );
   gpc1_1 gpc1_1_3116(
      {stage093[86]},
      {stage093[167]}
   );
   gpc1_1 gpc1_1_3117(
      {stage093[87]},
      {stage093[168]}
   );
   gpc1_1 gpc1_1_3118(
      {stage093[88]},
      {stage093[169]}
   );
   gpc1_1 gpc1_1_3119(
      {stage093[89]},
      {stage093[170]}
   );
   gpc1_1 gpc1_1_3120(
      {stage093[90]},
      {stage093[171]}
   );
   gpc1_1 gpc1_1_3121(
      {stage093[91]},
      {stage093[172]}
   );
   gpc1_1 gpc1_1_3122(
      {stage093[92]},
      {stage093[173]}
   );
   gpc1_1 gpc1_1_3123(
      {stage093[93]},
      {stage093[174]}
   );
   gpc1_1 gpc1_1_3124(
      {stage093[94]},
      {stage093[175]}
   );
   gpc1_1 gpc1_1_3125(
      {stage093[95]},
      {stage093[176]}
   );
   gpc1_1 gpc1_1_3126(
      {stage093[96]},
      {stage093[177]}
   );
   gpc1_1 gpc1_1_3127(
      {stage093[97]},
      {stage093[178]}
   );
   gpc1_1 gpc1_1_3128(
      {stage093[98]},
      {stage093[179]}
   );
   gpc1_1 gpc1_1_3129(
      {stage093[99]},
      {stage093[180]}
   );
   gpc1_1 gpc1_1_3130(
      {stage093[100]},
      {stage093[181]}
   );
   gpc1_1 gpc1_1_3131(
      {stage093[101]},
      {stage093[182]}
   );
   gpc1_1 gpc1_1_3132(
      {stage093[102]},
      {stage093[183]}
   );
   gpc1_1 gpc1_1_3133(
      {stage093[103]},
      {stage093[184]}
   );
   gpc606_5 gpc606_5_3134(
      {stage093[104], stage093[105], stage093[106], stage093[107], stage093[108], stage093[109]},
      {stage095[0], stage095[1], stage095[2], stage095[3], stage095[4], stage095[5]},
      {stage097[128], stage096[135], stage095[148], stage094[159], stage093[185]}
   );
   gpc606_5 gpc606_5_3135(
      {stage093[110], stage093[111], stage093[112], stage093[113], stage093[114], stage093[115]},
      {stage095[6], stage095[7], stage095[8], stage095[9], stage095[10], stage095[11]},
      {stage097[129], stage096[136], stage095[149], stage094[160], stage093[186]}
   );
   gpc606_5 gpc606_5_3136(
      {stage093[116], stage093[117], stage093[118], stage093[119], stage093[120], stage093[121]},
      {stage095[12], stage095[13], stage095[14], stage095[15], stage095[16], stage095[17]},
      {stage097[130], stage096[137], stage095[150], stage094[161], stage093[187]}
   );
   gpc606_5 gpc606_5_3137(
      {stage093[122], stage093[123], stage093[124], stage093[125], stage093[126], stage093[127]},
      {stage095[18], stage095[19], stage095[20], stage095[21], stage095[22], stage095[23]},
      {stage097[131], stage096[138], stage095[151], stage094[162], stage093[188]}
   );
   gpc1_1 gpc1_1_3138(
      {stage094[42]},
      {stage094[163]}
   );
   gpc1_1 gpc1_1_3139(
      {stage094[43]},
      {stage094[164]}
   );
   gpc1_1 gpc1_1_3140(
      {stage094[44]},
      {stage094[165]}
   );
   gpc1_1 gpc1_1_3141(
      {stage094[45]},
      {stage094[166]}
   );
   gpc1_1 gpc1_1_3142(
      {stage094[46]},
      {stage094[167]}
   );
   gpc1_1 gpc1_1_3143(
      {stage094[47]},
      {stage094[168]}
   );
   gpc1_1 gpc1_1_3144(
      {stage094[48]},
      {stage094[169]}
   );
   gpc1_1 gpc1_1_3145(
      {stage094[49]},
      {stage094[170]}
   );
   gpc1_1 gpc1_1_3146(
      {stage094[50]},
      {stage094[171]}
   );
   gpc1_1 gpc1_1_3147(
      {stage094[51]},
      {stage094[172]}
   );
   gpc1_1 gpc1_1_3148(
      {stage094[52]},
      {stage094[173]}
   );
   gpc1_1 gpc1_1_3149(
      {stage094[53]},
      {stage094[174]}
   );
   gpc1_1 gpc1_1_3150(
      {stage094[54]},
      {stage094[175]}
   );
   gpc1_1 gpc1_1_3151(
      {stage094[55]},
      {stage094[176]}
   );
   gpc1_1 gpc1_1_3152(
      {stage094[56]},
      {stage094[177]}
   );
   gpc1_1 gpc1_1_3153(
      {stage094[57]},
      {stage094[178]}
   );
   gpc1_1 gpc1_1_3154(
      {stage094[58]},
      {stage094[179]}
   );
   gpc1_1 gpc1_1_3155(
      {stage094[59]},
      {stage094[180]}
   );
   gpc1_1 gpc1_1_3156(
      {stage094[60]},
      {stage094[181]}
   );
   gpc1_1 gpc1_1_3157(
      {stage094[61]},
      {stage094[182]}
   );
   gpc1_1 gpc1_1_3158(
      {stage094[62]},
      {stage094[183]}
   );
   gpc606_5 gpc606_5_3159(
      {stage094[63], stage094[64], stage094[65], stage094[66], stage094[67], stage094[68]},
      {stage096[0], stage096[1], stage096[2], stage096[3], stage096[4], stage096[5]},
      {stage098[128], stage097[132], stage096[139], stage095[152], stage094[184]}
   );
   gpc606_5 gpc606_5_3160(
      {stage094[69], stage094[70], stage094[71], stage094[72], stage094[73], stage094[74]},
      {stage096[6], stage096[7], stage096[8], stage096[9], stage096[10], stage096[11]},
      {stage098[129], stage097[133], stage096[140], stage095[153], stage094[185]}
   );
   gpc606_5 gpc606_5_3161(
      {stage094[75], stage094[76], stage094[77], stage094[78], stage094[79], stage094[80]},
      {stage096[12], stage096[13], stage096[14], stage096[15], stage096[16], stage096[17]},
      {stage098[130], stage097[134], stage096[141], stage095[154], stage094[186]}
   );
   gpc606_5 gpc606_5_3162(
      {stage094[81], stage094[82], stage094[83], stage094[84], stage094[85], stage094[86]},
      {stage096[18], stage096[19], stage096[20], stage096[21], stage096[22], stage096[23]},
      {stage098[131], stage097[135], stage096[142], stage095[155], stage094[187]}
   );
   gpc606_5 gpc606_5_3163(
      {stage094[87], stage094[88], stage094[89], stage094[90], stage094[91], stage094[92]},
      {stage096[24], stage096[25], stage096[26], stage096[27], stage096[28], stage096[29]},
      {stage098[132], stage097[136], stage096[143], stage095[156], stage094[188]}
   );
   gpc606_5 gpc606_5_3164(
      {stage094[93], stage094[94], stage094[95], stage094[96], stage094[97], stage094[98]},
      {stage096[30], stage096[31], stage096[32], stage096[33], stage096[34], stage096[35]},
      {stage098[133], stage097[137], stage096[144], stage095[157], stage094[189]}
   );
   gpc606_5 gpc606_5_3165(
      {stage094[99], stage094[100], stage094[101], stage094[102], stage094[103], stage094[104]},
      {stage096[36], stage096[37], stage096[38], stage096[39], stage096[40], stage096[41]},
      {stage098[134], stage097[138], stage096[145], stage095[158], stage094[190]}
   );
   gpc606_5 gpc606_5_3166(
      {stage094[105], stage094[106], stage094[107], stage094[108], stage094[109], stage094[110]},
      {stage096[42], stage096[43], stage096[44], stage096[45], stage096[46], stage096[47]},
      {stage098[135], stage097[139], stage096[146], stage095[159], stage094[191]}
   );
   gpc606_5 gpc606_5_3167(
      {stage094[111], stage094[112], stage094[113], stage094[114], stage094[115], stage094[116]},
      {stage096[48], stage096[49], stage096[50], stage096[51], stage096[52], stage096[53]},
      {stage098[136], stage097[140], stage096[147], stage095[160], stage094[192]}
   );
   gpc606_5 gpc606_5_3168(
      {stage094[117], stage094[118], stage094[119], stage094[120], stage094[121], stage094[122]},
      {stage096[54], stage096[55], stage096[56], stage096[57], stage096[58], stage096[59]},
      {stage098[137], stage097[141], stage096[148], stage095[161], stage094[193]}
   );
   gpc615_5 gpc615_5_3169(
      {stage094[123], stage094[124], stage094[125], stage094[126], stage094[127]},
      {stage095[24]},
      {stage096[60], stage096[61], stage096[62], stage096[63], stage096[64], stage096[65]},
      {stage098[138], stage097[142], stage096[149], stage095[162], stage094[194]}
   );
   gpc1_1 gpc1_1_3170(
      {stage095[25]},
      {stage095[163]}
   );
   gpc606_5 gpc606_5_3171(
      {stage095[26], stage095[27], stage095[28], stage095[29], stage095[30], stage095[31]},
      {stage097[0], stage097[1], stage097[2], stage097[3], stage097[4], stage097[5]},
      {stage099[128], stage098[139], stage097[143], stage096[150], stage095[164]}
   );
   gpc606_5 gpc606_5_3172(
      {stage095[32], stage095[33], stage095[34], stage095[35], stage095[36], stage095[37]},
      {stage097[6], stage097[7], stage097[8], stage097[9], stage097[10], stage097[11]},
      {stage099[129], stage098[140], stage097[144], stage096[151], stage095[165]}
   );
   gpc606_5 gpc606_5_3173(
      {stage095[38], stage095[39], stage095[40], stage095[41], stage095[42], stage095[43]},
      {stage097[12], stage097[13], stage097[14], stage097[15], stage097[16], stage097[17]},
      {stage099[130], stage098[141], stage097[145], stage096[152], stage095[166]}
   );
   gpc606_5 gpc606_5_3174(
      {stage095[44], stage095[45], stage095[46], stage095[47], stage095[48], stage095[49]},
      {stage097[18], stage097[19], stage097[20], stage097[21], stage097[22], stage097[23]},
      {stage099[131], stage098[142], stage097[146], stage096[153], stage095[167]}
   );
   gpc606_5 gpc606_5_3175(
      {stage095[50], stage095[51], stage095[52], stage095[53], stage095[54], stage095[55]},
      {stage097[24], stage097[25], stage097[26], stage097[27], stage097[28], stage097[29]},
      {stage099[132], stage098[143], stage097[147], stage096[154], stage095[168]}
   );
   gpc606_5 gpc606_5_3176(
      {stage095[56], stage095[57], stage095[58], stage095[59], stage095[60], stage095[61]},
      {stage097[30], stage097[31], stage097[32], stage097[33], stage097[34], stage097[35]},
      {stage099[133], stage098[144], stage097[148], stage096[155], stage095[169]}
   );
   gpc606_5 gpc606_5_3177(
      {stage095[62], stage095[63], stage095[64], stage095[65], stage095[66], stage095[67]},
      {stage097[36], stage097[37], stage097[38], stage097[39], stage097[40], stage097[41]},
      {stage099[134], stage098[145], stage097[149], stage096[156], stage095[170]}
   );
   gpc606_5 gpc606_5_3178(
      {stage095[68], stage095[69], stage095[70], stage095[71], stage095[72], stage095[73]},
      {stage097[42], stage097[43], stage097[44], stage097[45], stage097[46], stage097[47]},
      {stage099[135], stage098[146], stage097[150], stage096[157], stage095[171]}
   );
   gpc606_5 gpc606_5_3179(
      {stage095[74], stage095[75], stage095[76], stage095[77], stage095[78], stage095[79]},
      {stage097[48], stage097[49], stage097[50], stage097[51], stage097[52], stage097[53]},
      {stage099[136], stage098[147], stage097[151], stage096[158], stage095[172]}
   );
   gpc606_5 gpc606_5_3180(
      {stage095[80], stage095[81], stage095[82], stage095[83], stage095[84], stage095[85]},
      {stage097[54], stage097[55], stage097[56], stage097[57], stage097[58], stage097[59]},
      {stage099[137], stage098[148], stage097[152], stage096[159], stage095[173]}
   );
   gpc606_5 gpc606_5_3181(
      {stage095[86], stage095[87], stage095[88], stage095[89], stage095[90], stage095[91]},
      {stage097[60], stage097[61], stage097[62], stage097[63], stage097[64], stage097[65]},
      {stage099[138], stage098[149], stage097[153], stage096[160], stage095[174]}
   );
   gpc606_5 gpc606_5_3182(
      {stage095[92], stage095[93], stage095[94], stage095[95], stage095[96], stage095[97]},
      {stage097[66], stage097[67], stage097[68], stage097[69], stage097[70], stage097[71]},
      {stage099[139], stage098[150], stage097[154], stage096[161], stage095[175]}
   );
   gpc606_5 gpc606_5_3183(
      {stage095[98], stage095[99], stage095[100], stage095[101], stage095[102], stage095[103]},
      {stage097[72], stage097[73], stage097[74], stage097[75], stage097[76], stage097[77]},
      {stage099[140], stage098[151], stage097[155], stage096[162], stage095[176]}
   );
   gpc606_5 gpc606_5_3184(
      {stage095[104], stage095[105], stage095[106], stage095[107], stage095[108], stage095[109]},
      {stage097[78], stage097[79], stage097[80], stage097[81], stage097[82], stage097[83]},
      {stage099[141], stage098[152], stage097[156], stage096[163], stage095[177]}
   );
   gpc606_5 gpc606_5_3185(
      {stage095[110], stage095[111], stage095[112], stage095[113], stage095[114], stage095[115]},
      {stage097[84], stage097[85], stage097[86], stage097[87], stage097[88], stage097[89]},
      {stage099[142], stage098[153], stage097[157], stage096[164], stage095[178]}
   );
   gpc606_5 gpc606_5_3186(
      {stage095[116], stage095[117], stage095[118], stage095[119], stage095[120], stage095[121]},
      {stage097[90], stage097[91], stage097[92], stage097[93], stage097[94], stage097[95]},
      {stage099[143], stage098[154], stage097[158], stage096[165], stage095[179]}
   );
   gpc606_5 gpc606_5_3187(
      {stage095[122], stage095[123], stage095[124], stage095[125], stage095[126], stage095[127]},
      {stage097[96], stage097[97], stage097[98], stage097[99], stage097[100], stage097[101]},
      {stage099[144], stage098[155], stage097[159], stage096[166], stage095[180]}
   );
   gpc1_1 gpc1_1_3188(
      {stage096[66]},
      {stage096[167]}
   );
   gpc1_1 gpc1_1_3189(
      {stage096[67]},
      {stage096[168]}
   );
   gpc1_1 gpc1_1_3190(
      {stage096[68]},
      {stage096[169]}
   );
   gpc1_1 gpc1_1_3191(
      {stage096[69]},
      {stage096[170]}
   );
   gpc1_1 gpc1_1_3192(
      {stage096[70]},
      {stage096[171]}
   );
   gpc1_1 gpc1_1_3193(
      {stage096[71]},
      {stage096[172]}
   );
   gpc1_1 gpc1_1_3194(
      {stage096[72]},
      {stage096[173]}
   );
   gpc1_1 gpc1_1_3195(
      {stage096[73]},
      {stage096[174]}
   );
   gpc606_5 gpc606_5_3196(
      {stage096[74], stage096[75], stage096[76], stage096[77], stage096[78], stage096[79]},
      {stage098[0], stage098[1], stage098[2], stage098[3], stage098[4], stage098[5]},
      {stage100[128], stage099[145], stage098[156], stage097[160], stage096[175]}
   );
   gpc606_5 gpc606_5_3197(
      {stage096[80], stage096[81], stage096[82], stage096[83], stage096[84], stage096[85]},
      {stage098[6], stage098[7], stage098[8], stage098[9], stage098[10], stage098[11]},
      {stage100[129], stage099[146], stage098[157], stage097[161], stage096[176]}
   );
   gpc606_5 gpc606_5_3198(
      {stage096[86], stage096[87], stage096[88], stage096[89], stage096[90], stage096[91]},
      {stage098[12], stage098[13], stage098[14], stage098[15], stage098[16], stage098[17]},
      {stage100[130], stage099[147], stage098[158], stage097[162], stage096[177]}
   );
   gpc606_5 gpc606_5_3199(
      {stage096[92], stage096[93], stage096[94], stage096[95], stage096[96], stage096[97]},
      {stage098[18], stage098[19], stage098[20], stage098[21], stage098[22], stage098[23]},
      {stage100[131], stage099[148], stage098[159], stage097[163], stage096[178]}
   );
   gpc606_5 gpc606_5_3200(
      {stage096[98], stage096[99], stage096[100], stage096[101], stage096[102], stage096[103]},
      {stage098[24], stage098[25], stage098[26], stage098[27], stage098[28], stage098[29]},
      {stage100[132], stage099[149], stage098[160], stage097[164], stage096[179]}
   );
   gpc606_5 gpc606_5_3201(
      {stage096[104], stage096[105], stage096[106], stage096[107], stage096[108], stage096[109]},
      {stage098[30], stage098[31], stage098[32], stage098[33], stage098[34], stage098[35]},
      {stage100[133], stage099[150], stage098[161], stage097[165], stage096[180]}
   );
   gpc606_5 gpc606_5_3202(
      {stage096[110], stage096[111], stage096[112], stage096[113], stage096[114], stage096[115]},
      {stage098[36], stage098[37], stage098[38], stage098[39], stage098[40], stage098[41]},
      {stage100[134], stage099[151], stage098[162], stage097[166], stage096[181]}
   );
   gpc606_5 gpc606_5_3203(
      {stage096[116], stage096[117], stage096[118], stage096[119], stage096[120], stage096[121]},
      {stage098[42], stage098[43], stage098[44], stage098[45], stage098[46], stage098[47]},
      {stage100[135], stage099[152], stage098[163], stage097[167], stage096[182]}
   );
   gpc606_5 gpc606_5_3204(
      {stage096[122], stage096[123], stage096[124], stage096[125], stage096[126], stage096[127]},
      {stage098[48], stage098[49], stage098[50], stage098[51], stage098[52], stage098[53]},
      {stage100[136], stage099[153], stage098[164], stage097[168], stage096[183]}
   );
   gpc1_1 gpc1_1_3205(
      {stage097[102]},
      {stage097[169]}
   );
   gpc615_5 gpc615_5_3206(
      {stage097[103], stage097[104], stage097[105], stage097[106], stage097[107]},
      {stage098[54]},
      {stage099[0], stage099[1], stage099[2], stage099[3], stage099[4], stage099[5]},
      {stage101[128], stage100[137], stage099[154], stage098[165], stage097[170]}
   );
   gpc615_5 gpc615_5_3207(
      {stage097[108], stage097[109], stage097[110], stage097[111], stage097[112]},
      {stage098[55]},
      {stage099[6], stage099[7], stage099[8], stage099[9], stage099[10], stage099[11]},
      {stage101[129], stage100[138], stage099[155], stage098[166], stage097[171]}
   );
   gpc615_5 gpc615_5_3208(
      {stage097[113], stage097[114], stage097[115], stage097[116], stage097[117]},
      {stage098[56]},
      {stage099[12], stage099[13], stage099[14], stage099[15], stage099[16], stage099[17]},
      {stage101[130], stage100[139], stage099[156], stage098[167], stage097[172]}
   );
   gpc615_5 gpc615_5_3209(
      {stage097[118], stage097[119], stage097[120], stage097[121], stage097[122]},
      {stage098[57]},
      {stage099[18], stage099[19], stage099[20], stage099[21], stage099[22], stage099[23]},
      {stage101[131], stage100[140], stage099[157], stage098[168], stage097[173]}
   );
   gpc615_5 gpc615_5_3210(
      {stage097[123], stage097[124], stage097[125], stage097[126], stage097[127]},
      {stage098[58]},
      {stage099[24], stage099[25], stage099[26], stage099[27], stage099[28], stage099[29]},
      {stage101[132], stage100[141], stage099[158], stage098[169], stage097[174]}
   );
   gpc1_1 gpc1_1_3211(
      {stage098[59]},
      {stage098[170]}
   );
   gpc1_1 gpc1_1_3212(
      {stage098[60]},
      {stage098[171]}
   );
   gpc1_1 gpc1_1_3213(
      {stage098[61]},
      {stage098[172]}
   );
   gpc606_5 gpc606_5_3214(
      {stage098[62], stage098[63], stage098[64], stage098[65], stage098[66], stage098[67]},
      {stage100[0], stage100[1], stage100[2], stage100[3], stage100[4], stage100[5]},
      {stage102[128], stage101[133], stage100[142], stage099[159], stage098[173]}
   );
   gpc606_5 gpc606_5_3215(
      {stage098[68], stage098[69], stage098[70], stage098[71], stage098[72], stage098[73]},
      {stage100[6], stage100[7], stage100[8], stage100[9], stage100[10], stage100[11]},
      {stage102[129], stage101[134], stage100[143], stage099[160], stage098[174]}
   );
   gpc606_5 gpc606_5_3216(
      {stage098[74], stage098[75], stage098[76], stage098[77], stage098[78], stage098[79]},
      {stage100[12], stage100[13], stage100[14], stage100[15], stage100[16], stage100[17]},
      {stage102[130], stage101[135], stage100[144], stage099[161], stage098[175]}
   );
   gpc606_5 gpc606_5_3217(
      {stage098[80], stage098[81], stage098[82], stage098[83], stage098[84], stage098[85]},
      {stage100[18], stage100[19], stage100[20], stage100[21], stage100[22], stage100[23]},
      {stage102[131], stage101[136], stage100[145], stage099[162], stage098[176]}
   );
   gpc606_5 gpc606_5_3218(
      {stage098[86], stage098[87], stage098[88], stage098[89], stage098[90], stage098[91]},
      {stage100[24], stage100[25], stage100[26], stage100[27], stage100[28], stage100[29]},
      {stage102[132], stage101[137], stage100[146], stage099[163], stage098[177]}
   );
   gpc606_5 gpc606_5_3219(
      {stage098[92], stage098[93], stage098[94], stage098[95], stage098[96], stage098[97]},
      {stage100[30], stage100[31], stage100[32], stage100[33], stage100[34], stage100[35]},
      {stage102[133], stage101[138], stage100[147], stage099[164], stage098[178]}
   );
   gpc606_5 gpc606_5_3220(
      {stage098[98], stage098[99], stage098[100], stage098[101], stage098[102], stage098[103]},
      {stage100[36], stage100[37], stage100[38], stage100[39], stage100[40], stage100[41]},
      {stage102[134], stage101[139], stage100[148], stage099[165], stage098[179]}
   );
   gpc606_5 gpc606_5_3221(
      {stage098[104], stage098[105], stage098[106], stage098[107], stage098[108], stage098[109]},
      {stage100[42], stage100[43], stage100[44], stage100[45], stage100[46], stage100[47]},
      {stage102[135], stage101[140], stage100[149], stage099[166], stage098[180]}
   );
   gpc606_5 gpc606_5_3222(
      {stage098[110], stage098[111], stage098[112], stage098[113], stage098[114], stage098[115]},
      {stage100[48], stage100[49], stage100[50], stage100[51], stage100[52], stage100[53]},
      {stage102[136], stage101[141], stage100[150], stage099[167], stage098[181]}
   );
   gpc606_5 gpc606_5_3223(
      {stage098[116], stage098[117], stage098[118], stage098[119], stage098[120], stage098[121]},
      {stage100[54], stage100[55], stage100[56], stage100[57], stage100[58], stage100[59]},
      {stage102[137], stage101[142], stage100[151], stage099[168], stage098[182]}
   );
   gpc606_5 gpc606_5_3224(
      {stage098[122], stage098[123], stage098[124], stage098[125], stage098[126], stage098[127]},
      {stage100[60], stage100[61], stage100[62], stage100[63], stage100[64], stage100[65]},
      {stage102[138], stage101[143], stage100[152], stage099[169], stage098[183]}
   );
   gpc1_1 gpc1_1_3225(
      {stage099[30]},
      {stage099[170]}
   );
   gpc1_1 gpc1_1_3226(
      {stage099[31]},
      {stage099[171]}
   );
   gpc1_1 gpc1_1_3227(
      {stage099[32]},
      {stage099[172]}
   );
   gpc1_1 gpc1_1_3228(
      {stage099[33]},
      {stage099[173]}
   );
   gpc1_1 gpc1_1_3229(
      {stage099[34]},
      {stage099[174]}
   );
   gpc1_1 gpc1_1_3230(
      {stage099[35]},
      {stage099[175]}
   );
   gpc1_1 gpc1_1_3231(
      {stage099[36]},
      {stage099[176]}
   );
   gpc1_1 gpc1_1_3232(
      {stage099[37]},
      {stage099[177]}
   );
   gpc1_1 gpc1_1_3233(
      {stage099[38]},
      {stage099[178]}
   );
   gpc1_1 gpc1_1_3234(
      {stage099[39]},
      {stage099[179]}
   );
   gpc1_1 gpc1_1_3235(
      {stage099[40]},
      {stage099[180]}
   );
   gpc1_1 gpc1_1_3236(
      {stage099[41]},
      {stage099[181]}
   );
   gpc1_1 gpc1_1_3237(
      {stage099[42]},
      {stage099[182]}
   );
   gpc1_1 gpc1_1_3238(
      {stage099[43]},
      {stage099[183]}
   );
   gpc1_1 gpc1_1_3239(
      {stage099[44]},
      {stage099[184]}
   );
   gpc1_1 gpc1_1_3240(
      {stage099[45]},
      {stage099[185]}
   );
   gpc1_1 gpc1_1_3241(
      {stage099[46]},
      {stage099[186]}
   );
   gpc1_1 gpc1_1_3242(
      {stage099[47]},
      {stage099[187]}
   );
   gpc1_1 gpc1_1_3243(
      {stage099[48]},
      {stage099[188]}
   );
   gpc1_1 gpc1_1_3244(
      {stage099[49]},
      {stage099[189]}
   );
   gpc1_1 gpc1_1_3245(
      {stage099[50]},
      {stage099[190]}
   );
   gpc606_5 gpc606_5_3246(
      {stage099[51], stage099[52], stage099[53], stage099[54], stage099[55], stage099[56]},
      {stage101[0], stage101[1], stage101[2], stage101[3], stage101[4], stage101[5]},
      {stage103[128], stage102[139], stage101[144], stage100[153], stage099[191]}
   );
   gpc606_5 gpc606_5_3247(
      {stage099[57], stage099[58], stage099[59], stage099[60], stage099[61], stage099[62]},
      {stage101[6], stage101[7], stage101[8], stage101[9], stage101[10], stage101[11]},
      {stage103[129], stage102[140], stage101[145], stage100[154], stage099[192]}
   );
   gpc606_5 gpc606_5_3248(
      {stage099[63], stage099[64], stage099[65], stage099[66], stage099[67], stage099[68]},
      {stage101[12], stage101[13], stage101[14], stage101[15], stage101[16], stage101[17]},
      {stage103[130], stage102[141], stage101[146], stage100[155], stage099[193]}
   );
   gpc606_5 gpc606_5_3249(
      {stage099[69], stage099[70], stage099[71], stage099[72], stage099[73], stage099[74]},
      {stage101[18], stage101[19], stage101[20], stage101[21], stage101[22], stage101[23]},
      {stage103[131], stage102[142], stage101[147], stage100[156], stage099[194]}
   );
   gpc606_5 gpc606_5_3250(
      {stage099[75], stage099[76], stage099[77], stage099[78], stage099[79], stage099[80]},
      {stage101[24], stage101[25], stage101[26], stage101[27], stage101[28], stage101[29]},
      {stage103[132], stage102[143], stage101[148], stage100[157], stage099[195]}
   );
   gpc606_5 gpc606_5_3251(
      {stage099[81], stage099[82], stage099[83], stage099[84], stage099[85], stage099[86]},
      {stage101[30], stage101[31], stage101[32], stage101[33], stage101[34], stage101[35]},
      {stage103[133], stage102[144], stage101[149], stage100[158], stage099[196]}
   );
   gpc606_5 gpc606_5_3252(
      {stage099[87], stage099[88], stage099[89], stage099[90], stage099[91], stage099[92]},
      {stage101[36], stage101[37], stage101[38], stage101[39], stage101[40], stage101[41]},
      {stage103[134], stage102[145], stage101[150], stage100[159], stage099[197]}
   );
   gpc606_5 gpc606_5_3253(
      {stage099[93], stage099[94], stage099[95], stage099[96], stage099[97], stage099[98]},
      {stage101[42], stage101[43], stage101[44], stage101[45], stage101[46], stage101[47]},
      {stage103[135], stage102[146], stage101[151], stage100[160], stage099[198]}
   );
   gpc606_5 gpc606_5_3254(
      {stage099[99], stage099[100], stage099[101], stage099[102], stage099[103], stage099[104]},
      {stage101[48], stage101[49], stage101[50], stage101[51], stage101[52], stage101[53]},
      {stage103[136], stage102[147], stage101[152], stage100[161], stage099[199]}
   );
   gpc606_5 gpc606_5_3255(
      {stage099[105], stage099[106], stage099[107], stage099[108], stage099[109], stage099[110]},
      {stage101[54], stage101[55], stage101[56], stage101[57], stage101[58], stage101[59]},
      {stage103[137], stage102[148], stage101[153], stage100[162], stage099[200]}
   );
   gpc606_5 gpc606_5_3256(
      {stage099[111], stage099[112], stage099[113], stage099[114], stage099[115], stage099[116]},
      {stage101[60], stage101[61], stage101[62], stage101[63], stage101[64], stage101[65]},
      {stage103[138], stage102[149], stage101[154], stage100[163], stage099[201]}
   );
   gpc606_5 gpc606_5_3257(
      {stage099[117], stage099[118], stage099[119], stage099[120], stage099[121], stage099[122]},
      {stage101[66], stage101[67], stage101[68], stage101[69], stage101[70], stage101[71]},
      {stage103[139], stage102[150], stage101[155], stage100[164], stage099[202]}
   );
   gpc615_5 gpc615_5_3258(
      {stage099[123], stage099[124], stage099[125], stage099[126], stage099[127]},
      {stage100[66]},
      {stage101[72], stage101[73], stage101[74], stage101[75], stage101[76], stage101[77]},
      {stage103[140], stage102[151], stage101[156], stage100[165], stage099[203]}
   );
   gpc1_1 gpc1_1_3259(
      {stage100[67]},
      {stage100[166]}
   );
   gpc606_5 gpc606_5_3260(
      {stage100[68], stage100[69], stage100[70], stage100[71], stage100[72], stage100[73]},
      {stage102[0], stage102[1], stage102[2], stage102[3], stage102[4], stage102[5]},
      {stage104[128], stage103[141], stage102[152], stage101[157], stage100[167]}
   );
   gpc606_5 gpc606_5_3261(
      {stage100[74], stage100[75], stage100[76], stage100[77], stage100[78], stage100[79]},
      {stage102[6], stage102[7], stage102[8], stage102[9], stage102[10], stage102[11]},
      {stage104[129], stage103[142], stage102[153], stage101[158], stage100[168]}
   );
   gpc606_5 gpc606_5_3262(
      {stage100[80], stage100[81], stage100[82], stage100[83], stage100[84], stage100[85]},
      {stage102[12], stage102[13], stage102[14], stage102[15], stage102[16], stage102[17]},
      {stage104[130], stage103[143], stage102[154], stage101[159], stage100[169]}
   );
   gpc606_5 gpc606_5_3263(
      {stage100[86], stage100[87], stage100[88], stage100[89], stage100[90], stage100[91]},
      {stage102[18], stage102[19], stage102[20], stage102[21], stage102[22], stage102[23]},
      {stage104[131], stage103[144], stage102[155], stage101[160], stage100[170]}
   );
   gpc606_5 gpc606_5_3264(
      {stage100[92], stage100[93], stage100[94], stage100[95], stage100[96], stage100[97]},
      {stage102[24], stage102[25], stage102[26], stage102[27], stage102[28], stage102[29]},
      {stage104[132], stage103[145], stage102[156], stage101[161], stage100[171]}
   );
   gpc615_5 gpc615_5_3265(
      {stage100[98], stage100[99], stage100[100], stage100[101], stage100[102]},
      {stage101[78]},
      {stage102[30], stage102[31], stage102[32], stage102[33], stage102[34], stage102[35]},
      {stage104[133], stage103[146], stage102[157], stage101[162], stage100[172]}
   );
   gpc615_5 gpc615_5_3266(
      {stage100[103], stage100[104], stage100[105], stage100[106], stage100[107]},
      {stage101[79]},
      {stage102[36], stage102[37], stage102[38], stage102[39], stage102[40], stage102[41]},
      {stage104[134], stage103[147], stage102[158], stage101[163], stage100[173]}
   );
   gpc615_5 gpc615_5_3267(
      {stage100[108], stage100[109], stage100[110], stage100[111], stage100[112]},
      {stage101[80]},
      {stage102[42], stage102[43], stage102[44], stage102[45], stage102[46], stage102[47]},
      {stage104[135], stage103[148], stage102[159], stage101[164], stage100[174]}
   );
   gpc615_5 gpc615_5_3268(
      {stage100[113], stage100[114], stage100[115], stage100[116], stage100[117]},
      {stage101[81]},
      {stage102[48], stage102[49], stage102[50], stage102[51], stage102[52], stage102[53]},
      {stage104[136], stage103[149], stage102[160], stage101[165], stage100[175]}
   );
   gpc615_5 gpc615_5_3269(
      {stage100[118], stage100[119], stage100[120], stage100[121], stage100[122]},
      {stage101[82]},
      {stage102[54], stage102[55], stage102[56], stage102[57], stage102[58], stage102[59]},
      {stage104[137], stage103[150], stage102[161], stage101[166], stage100[176]}
   );
   gpc615_5 gpc615_5_3270(
      {stage100[123], stage100[124], stage100[125], stage100[126], stage100[127]},
      {stage101[83]},
      {stage102[60], stage102[61], stage102[62], stage102[63], stage102[64], stage102[65]},
      {stage104[138], stage103[151], stage102[162], stage101[167], stage100[177]}
   );
   gpc1_1 gpc1_1_3271(
      {stage101[84]},
      {stage101[168]}
   );
   gpc1_1 gpc1_1_3272(
      {stage101[85]},
      {stage101[169]}
   );
   gpc1_1 gpc1_1_3273(
      {stage101[86]},
      {stage101[170]}
   );
   gpc1_1 gpc1_1_3274(
      {stage101[87]},
      {stage101[171]}
   );
   gpc1_1 gpc1_1_3275(
      {stage101[88]},
      {stage101[172]}
   );
   gpc1_1 gpc1_1_3276(
      {stage101[89]},
      {stage101[173]}
   );
   gpc1_1 gpc1_1_3277(
      {stage101[90]},
      {stage101[174]}
   );
   gpc1_1 gpc1_1_3278(
      {stage101[91]},
      {stage101[175]}
   );
   gpc1_1 gpc1_1_3279(
      {stage101[92]},
      {stage101[176]}
   );
   gpc1_1 gpc1_1_3280(
      {stage101[93]},
      {stage101[177]}
   );
   gpc1_1 gpc1_1_3281(
      {stage101[94]},
      {stage101[178]}
   );
   gpc1_1 gpc1_1_3282(
      {stage101[95]},
      {stage101[179]}
   );
   gpc1_1 gpc1_1_3283(
      {stage101[96]},
      {stage101[180]}
   );
   gpc1_1 gpc1_1_3284(
      {stage101[97]},
      {stage101[181]}
   );
   gpc1_1 gpc1_1_3285(
      {stage101[98]},
      {stage101[182]}
   );
   gpc1_1 gpc1_1_3286(
      {stage101[99]},
      {stage101[183]}
   );
   gpc1_1 gpc1_1_3287(
      {stage101[100]},
      {stage101[184]}
   );
   gpc1_1 gpc1_1_3288(
      {stage101[101]},
      {stage101[185]}
   );
   gpc1_1 gpc1_1_3289(
      {stage101[102]},
      {stage101[186]}
   );
   gpc1_1 gpc1_1_3290(
      {stage101[103]},
      {stage101[187]}
   );
   gpc606_5 gpc606_5_3291(
      {stage101[104], stage101[105], stage101[106], stage101[107], stage101[108], stage101[109]},
      {stage103[0], stage103[1], stage103[2], stage103[3], stage103[4], stage103[5]},
      {stage105[128], stage104[139], stage103[152], stage102[163], stage101[188]}
   );
   gpc606_5 gpc606_5_3292(
      {stage101[110], stage101[111], stage101[112], stage101[113], stage101[114], stage101[115]},
      {stage103[6], stage103[7], stage103[8], stage103[9], stage103[10], stage103[11]},
      {stage105[129], stage104[140], stage103[153], stage102[164], stage101[189]}
   );
   gpc606_5 gpc606_5_3293(
      {stage101[116], stage101[117], stage101[118], stage101[119], stage101[120], stage101[121]},
      {stage103[12], stage103[13], stage103[14], stage103[15], stage103[16], stage103[17]},
      {stage105[130], stage104[141], stage103[154], stage102[165], stage101[190]}
   );
   gpc606_5 gpc606_5_3294(
      {stage101[122], stage101[123], stage101[124], stage101[125], stage101[126], stage101[127]},
      {stage103[18], stage103[19], stage103[20], stage103[21], stage103[22], stage103[23]},
      {stage105[131], stage104[142], stage103[155], stage102[166], stage101[191]}
   );
   gpc1_1 gpc1_1_3295(
      {stage102[66]},
      {stage102[167]}
   );
   gpc1_1 gpc1_1_3296(
      {stage102[67]},
      {stage102[168]}
   );
   gpc1_1 gpc1_1_3297(
      {stage102[68]},
      {stage102[169]}
   );
   gpc1_1 gpc1_1_3298(
      {stage102[69]},
      {stage102[170]}
   );
   gpc1_1 gpc1_1_3299(
      {stage102[70]},
      {stage102[171]}
   );
   gpc1_1 gpc1_1_3300(
      {stage102[71]},
      {stage102[172]}
   );
   gpc1_1 gpc1_1_3301(
      {stage102[72]},
      {stage102[173]}
   );
   gpc1_1 gpc1_1_3302(
      {stage102[73]},
      {stage102[174]}
   );
   gpc1_1 gpc1_1_3303(
      {stage102[74]},
      {stage102[175]}
   );
   gpc1_1 gpc1_1_3304(
      {stage102[75]},
      {stage102[176]}
   );
   gpc1_1 gpc1_1_3305(
      {stage102[76]},
      {stage102[177]}
   );
   gpc1_1 gpc1_1_3306(
      {stage102[77]},
      {stage102[178]}
   );
   gpc1_1 gpc1_1_3307(
      {stage102[78]},
      {stage102[179]}
   );
   gpc1_1 gpc1_1_3308(
      {stage102[79]},
      {stage102[180]}
   );
   gpc1_1 gpc1_1_3309(
      {stage102[80]},
      {stage102[181]}
   );
   gpc1_1 gpc1_1_3310(
      {stage102[81]},
      {stage102[182]}
   );
   gpc1_1 gpc1_1_3311(
      {stage102[82]},
      {stage102[183]}
   );
   gpc1_1 gpc1_1_3312(
      {stage102[83]},
      {stage102[184]}
   );
   gpc1_1 gpc1_1_3313(
      {stage102[84]},
      {stage102[185]}
   );
   gpc1_1 gpc1_1_3314(
      {stage102[85]},
      {stage102[186]}
   );
   gpc1_1 gpc1_1_3315(
      {stage102[86]},
      {stage102[187]}
   );
   gpc1_1 gpc1_1_3316(
      {stage102[87]},
      {stage102[188]}
   );
   gpc1_1 gpc1_1_3317(
      {stage102[88]},
      {stage102[189]}
   );
   gpc1_1 gpc1_1_3318(
      {stage102[89]},
      {stage102[190]}
   );
   gpc1_1 gpc1_1_3319(
      {stage102[90]},
      {stage102[191]}
   );
   gpc1_1 gpc1_1_3320(
      {stage102[91]},
      {stage102[192]}
   );
   gpc1_1 gpc1_1_3321(
      {stage102[92]},
      {stage102[193]}
   );
   gpc606_5 gpc606_5_3322(
      {stage102[93], stage102[94], stage102[95], stage102[96], stage102[97], stage102[98]},
      {stage104[0], stage104[1], stage104[2], stage104[3], stage104[4], stage104[5]},
      {stage106[128], stage105[132], stage104[143], stage103[156], stage102[194]}
   );
   gpc606_5 gpc606_5_3323(
      {stage102[99], stage102[100], stage102[101], stage102[102], stage102[103], stage102[104]},
      {stage104[6], stage104[7], stage104[8], stage104[9], stage104[10], stage104[11]},
      {stage106[129], stage105[133], stage104[144], stage103[157], stage102[195]}
   );
   gpc606_5 gpc606_5_3324(
      {stage102[105], stage102[106], stage102[107], stage102[108], stage102[109], stage102[110]},
      {stage104[12], stage104[13], stage104[14], stage104[15], stage104[16], stage104[17]},
      {stage106[130], stage105[134], stage104[145], stage103[158], stage102[196]}
   );
   gpc606_5 gpc606_5_3325(
      {stage102[111], stage102[112], stage102[113], stage102[114], stage102[115], stage102[116]},
      {stage104[18], stage104[19], stage104[20], stage104[21], stage104[22], stage104[23]},
      {stage106[131], stage105[135], stage104[146], stage103[159], stage102[197]}
   );
   gpc606_5 gpc606_5_3326(
      {stage102[117], stage102[118], stage102[119], stage102[120], stage102[121], stage102[122]},
      {stage104[24], stage104[25], stage104[26], stage104[27], stage104[28], stage104[29]},
      {stage106[132], stage105[136], stage104[147], stage103[160], stage102[198]}
   );
   gpc615_5 gpc615_5_3327(
      {stage102[123], stage102[124], stage102[125], stage102[126], stage102[127]},
      {stage103[24]},
      {stage104[30], stage104[31], stage104[32], stage104[33], stage104[34], stage104[35]},
      {stage106[133], stage105[137], stage104[148], stage103[161], stage102[199]}
   );
   gpc1_1 gpc1_1_3328(
      {stage103[25]},
      {stage103[162]}
   );
   gpc1_1 gpc1_1_3329(
      {stage103[26]},
      {stage103[163]}
   );
   gpc1_1 gpc1_1_3330(
      {stage103[27]},
      {stage103[164]}
   );
   gpc1_1 gpc1_1_3331(
      {stage103[28]},
      {stage103[165]}
   );
   gpc1_1 gpc1_1_3332(
      {stage103[29]},
      {stage103[166]}
   );
   gpc1_1 gpc1_1_3333(
      {stage103[30]},
      {stage103[167]}
   );
   gpc1_1 gpc1_1_3334(
      {stage103[31]},
      {stage103[168]}
   );
   gpc1_1 gpc1_1_3335(
      {stage103[32]},
      {stage103[169]}
   );
   gpc1_1 gpc1_1_3336(
      {stage103[33]},
      {stage103[170]}
   );
   gpc1_1 gpc1_1_3337(
      {stage103[34]},
      {stage103[171]}
   );
   gpc1_1 gpc1_1_3338(
      {stage103[35]},
      {stage103[172]}
   );
   gpc1_1 gpc1_1_3339(
      {stage103[36]},
      {stage103[173]}
   );
   gpc1_1 gpc1_1_3340(
      {stage103[37]},
      {stage103[174]}
   );
   gpc606_5 gpc606_5_3341(
      {stage103[38], stage103[39], stage103[40], stage103[41], stage103[42], stage103[43]},
      {stage105[0], stage105[1], stage105[2], stage105[3], stage105[4], stage105[5]},
      {stage107[128], stage106[134], stage105[138], stage104[149], stage103[175]}
   );
   gpc606_5 gpc606_5_3342(
      {stage103[44], stage103[45], stage103[46], stage103[47], stage103[48], stage103[49]},
      {stage105[6], stage105[7], stage105[8], stage105[9], stage105[10], stage105[11]},
      {stage107[129], stage106[135], stage105[139], stage104[150], stage103[176]}
   );
   gpc606_5 gpc606_5_3343(
      {stage103[50], stage103[51], stage103[52], stage103[53], stage103[54], stage103[55]},
      {stage105[12], stage105[13], stage105[14], stage105[15], stage105[16], stage105[17]},
      {stage107[130], stage106[136], stage105[140], stage104[151], stage103[177]}
   );
   gpc606_5 gpc606_5_3344(
      {stage103[56], stage103[57], stage103[58], stage103[59], stage103[60], stage103[61]},
      {stage105[18], stage105[19], stage105[20], stage105[21], stage105[22], stage105[23]},
      {stage107[131], stage106[137], stage105[141], stage104[152], stage103[178]}
   );
   gpc606_5 gpc606_5_3345(
      {stage103[62], stage103[63], stage103[64], stage103[65], stage103[66], stage103[67]},
      {stage105[24], stage105[25], stage105[26], stage105[27], stage105[28], stage105[29]},
      {stage107[132], stage106[138], stage105[142], stage104[153], stage103[179]}
   );
   gpc615_5 gpc615_5_3346(
      {stage103[68], stage103[69], stage103[70], stage103[71], stage103[72]},
      {stage104[36]},
      {stage105[30], stage105[31], stage105[32], stage105[33], stage105[34], stage105[35]},
      {stage107[133], stage106[139], stage105[143], stage104[154], stage103[180]}
   );
   gpc615_5 gpc615_5_3347(
      {stage103[73], stage103[74], stage103[75], stage103[76], stage103[77]},
      {stage104[37]},
      {stage105[36], stage105[37], stage105[38], stage105[39], stage105[40], stage105[41]},
      {stage107[134], stage106[140], stage105[144], stage104[155], stage103[181]}
   );
   gpc615_5 gpc615_5_3348(
      {stage103[78], stage103[79], stage103[80], stage103[81], stage103[82]},
      {stage104[38]},
      {stage105[42], stage105[43], stage105[44], stage105[45], stage105[46], stage105[47]},
      {stage107[135], stage106[141], stage105[145], stage104[156], stage103[182]}
   );
   gpc615_5 gpc615_5_3349(
      {stage103[83], stage103[84], stage103[85], stage103[86], stage103[87]},
      {stage104[39]},
      {stage105[48], stage105[49], stage105[50], stage105[51], stage105[52], stage105[53]},
      {stage107[136], stage106[142], stage105[146], stage104[157], stage103[183]}
   );
   gpc615_5 gpc615_5_3350(
      {stage103[88], stage103[89], stage103[90], stage103[91], stage103[92]},
      {stage104[40]},
      {stage105[54], stage105[55], stage105[56], stage105[57], stage105[58], stage105[59]},
      {stage107[137], stage106[143], stage105[147], stage104[158], stage103[184]}
   );
   gpc615_5 gpc615_5_3351(
      {stage103[93], stage103[94], stage103[95], stage103[96], stage103[97]},
      {stage104[41]},
      {stage105[60], stage105[61], stage105[62], stage105[63], stage105[64], stage105[65]},
      {stage107[138], stage106[144], stage105[148], stage104[159], stage103[185]}
   );
   gpc615_5 gpc615_5_3352(
      {stage103[98], stage103[99], stage103[100], stage103[101], stage103[102]},
      {stage104[42]},
      {stage105[66], stage105[67], stage105[68], stage105[69], stage105[70], stage105[71]},
      {stage107[139], stage106[145], stage105[149], stage104[160], stage103[186]}
   );
   gpc615_5 gpc615_5_3353(
      {stage103[103], stage103[104], stage103[105], stage103[106], stage103[107]},
      {stage104[43]},
      {stage105[72], stage105[73], stage105[74], stage105[75], stage105[76], stage105[77]},
      {stage107[140], stage106[146], stage105[150], stage104[161], stage103[187]}
   );
   gpc615_5 gpc615_5_3354(
      {stage103[108], stage103[109], stage103[110], stage103[111], stage103[112]},
      {stage104[44]},
      {stage105[78], stage105[79], stage105[80], stage105[81], stage105[82], stage105[83]},
      {stage107[141], stage106[147], stage105[151], stage104[162], stage103[188]}
   );
   gpc615_5 gpc615_5_3355(
      {stage103[113], stage103[114], stage103[115], stage103[116], stage103[117]},
      {stage104[45]},
      {stage105[84], stage105[85], stage105[86], stage105[87], stage105[88], stage105[89]},
      {stage107[142], stage106[148], stage105[152], stage104[163], stage103[189]}
   );
   gpc615_5 gpc615_5_3356(
      {stage103[118], stage103[119], stage103[120], stage103[121], stage103[122]},
      {stage104[46]},
      {stage105[90], stage105[91], stage105[92], stage105[93], stage105[94], stage105[95]},
      {stage107[143], stage106[149], stage105[153], stage104[164], stage103[190]}
   );
   gpc615_5 gpc615_5_3357(
      {stage103[123], stage103[124], stage103[125], stage103[126], stage103[127]},
      {stage104[47]},
      {stage105[96], stage105[97], stage105[98], stage105[99], stage105[100], stage105[101]},
      {stage107[144], stage106[150], stage105[154], stage104[165], stage103[191]}
   );
   gpc1_1 gpc1_1_3358(
      {stage104[48]},
      {stage104[166]}
   );
   gpc1_1 gpc1_1_3359(
      {stage104[49]},
      {stage104[167]}
   );
   gpc1_1 gpc1_1_3360(
      {stage104[50]},
      {stage104[168]}
   );
   gpc1_1 gpc1_1_3361(
      {stage104[51]},
      {stage104[169]}
   );
   gpc1_1 gpc1_1_3362(
      {stage104[52]},
      {stage104[170]}
   );
   gpc1_1 gpc1_1_3363(
      {stage104[53]},
      {stage104[171]}
   );
   gpc1_1 gpc1_1_3364(
      {stage104[54]},
      {stage104[172]}
   );
   gpc1_1 gpc1_1_3365(
      {stage104[55]},
      {stage104[173]}
   );
   gpc1_1 gpc1_1_3366(
      {stage104[56]},
      {stage104[174]}
   );
   gpc1_1 gpc1_1_3367(
      {stage104[57]},
      {stage104[175]}
   );
   gpc1_1 gpc1_1_3368(
      {stage104[58]},
      {stage104[176]}
   );
   gpc1_1 gpc1_1_3369(
      {stage104[59]},
      {stage104[177]}
   );
   gpc1_1 gpc1_1_3370(
      {stage104[60]},
      {stage104[178]}
   );
   gpc1_1 gpc1_1_3371(
      {stage104[61]},
      {stage104[179]}
   );
   gpc1_1 gpc1_1_3372(
      {stage104[62]},
      {stage104[180]}
   );
   gpc1_1 gpc1_1_3373(
      {stage104[63]},
      {stage104[181]}
   );
   gpc1_1 gpc1_1_3374(
      {stage104[64]},
      {stage104[182]}
   );
   gpc1_1 gpc1_1_3375(
      {stage104[65]},
      {stage104[183]}
   );
   gpc1_1 gpc1_1_3376(
      {stage104[66]},
      {stage104[184]}
   );
   gpc1_1 gpc1_1_3377(
      {stage104[67]},
      {stage104[185]}
   );
   gpc1_1 gpc1_1_3378(
      {stage104[68]},
      {stage104[186]}
   );
   gpc1_1 gpc1_1_3379(
      {stage104[69]},
      {stage104[187]}
   );
   gpc1_1 gpc1_1_3380(
      {stage104[70]},
      {stage104[188]}
   );
   gpc1_1 gpc1_1_3381(
      {stage104[71]},
      {stage104[189]}
   );
   gpc1_1 gpc1_1_3382(
      {stage104[72]},
      {stage104[190]}
   );
   gpc1_1 gpc1_1_3383(
      {stage104[73]},
      {stage104[191]}
   );
   gpc1_1 gpc1_1_3384(
      {stage104[74]},
      {stage104[192]}
   );
   gpc1_1 gpc1_1_3385(
      {stage104[75]},
      {stage104[193]}
   );
   gpc1_1 gpc1_1_3386(
      {stage104[76]},
      {stage104[194]}
   );
   gpc1_1 gpc1_1_3387(
      {stage104[77]},
      {stage104[195]}
   );
   gpc1_1 gpc1_1_3388(
      {stage104[78]},
      {stage104[196]}
   );
   gpc1_1 gpc1_1_3389(
      {stage104[79]},
      {stage104[197]}
   );
   gpc1_1 gpc1_1_3390(
      {stage104[80]},
      {stage104[198]}
   );
   gpc1_1 gpc1_1_3391(
      {stage104[81]},
      {stage104[199]}
   );
   gpc1_1 gpc1_1_3392(
      {stage104[82]},
      {stage104[200]}
   );
   gpc1_1 gpc1_1_3393(
      {stage104[83]},
      {stage104[201]}
   );
   gpc1_1 gpc1_1_3394(
      {stage104[84]},
      {stage104[202]}
   );
   gpc1_1 gpc1_1_3395(
      {stage104[85]},
      {stage104[203]}
   );
   gpc606_5 gpc606_5_3396(
      {stage104[86], stage104[87], stage104[88], stage104[89], stage104[90], stage104[91]},
      {stage106[0], stage106[1], stage106[2], stage106[3], stage106[4], stage106[5]},
      {stage108[128], stage107[145], stage106[151], stage105[155], stage104[204]}
   );
   gpc606_5 gpc606_5_3397(
      {stage104[92], stage104[93], stage104[94], stage104[95], stage104[96], stage104[97]},
      {stage106[6], stage106[7], stage106[8], stage106[9], stage106[10], stage106[11]},
      {stage108[129], stage107[146], stage106[152], stage105[156], stage104[205]}
   );
   gpc606_5 gpc606_5_3398(
      {stage104[98], stage104[99], stage104[100], stage104[101], stage104[102], stage104[103]},
      {stage106[12], stage106[13], stage106[14], stage106[15], stage106[16], stage106[17]},
      {stage108[130], stage107[147], stage106[153], stage105[157], stage104[206]}
   );
   gpc606_5 gpc606_5_3399(
      {stage104[104], stage104[105], stage104[106], stage104[107], stage104[108], stage104[109]},
      {stage106[18], stage106[19], stage106[20], stage106[21], stage106[22], stage106[23]},
      {stage108[131], stage107[148], stage106[154], stage105[158], stage104[207]}
   );
   gpc606_5 gpc606_5_3400(
      {stage104[110], stage104[111], stage104[112], stage104[113], stage104[114], stage104[115]},
      {stage106[24], stage106[25], stage106[26], stage106[27], stage106[28], stage106[29]},
      {stage108[132], stage107[149], stage106[155], stage105[159], stage104[208]}
   );
   gpc606_5 gpc606_5_3401(
      {stage104[116], stage104[117], stage104[118], stage104[119], stage104[120], stage104[121]},
      {stage106[30], stage106[31], stage106[32], stage106[33], stage106[34], stage106[35]},
      {stage108[133], stage107[150], stage106[156], stage105[160], stage104[209]}
   );
   gpc606_5 gpc606_5_3402(
      {stage104[122], stage104[123], stage104[124], stage104[125], stage104[126], stage104[127]},
      {stage106[36], stage106[37], stage106[38], stage106[39], stage106[40], stage106[41]},
      {stage108[134], stage107[151], stage106[157], stage105[161], stage104[210]}
   );
   gpc1_1 gpc1_1_3403(
      {stage105[102]},
      {stage105[162]}
   );
   gpc1_1 gpc1_1_3404(
      {stage105[103]},
      {stage105[163]}
   );
   gpc1_1 gpc1_1_3405(
      {stage105[104]},
      {stage105[164]}
   );
   gpc1_1 gpc1_1_3406(
      {stage105[105]},
      {stage105[165]}
   );
   gpc1_1 gpc1_1_3407(
      {stage105[106]},
      {stage105[166]}
   );
   gpc1_1 gpc1_1_3408(
      {stage105[107]},
      {stage105[167]}
   );
   gpc1_1 gpc1_1_3409(
      {stage105[108]},
      {stage105[168]}
   );
   gpc1_1 gpc1_1_3410(
      {stage105[109]},
      {stage105[169]}
   );
   gpc1_1 gpc1_1_3411(
      {stage105[110]},
      {stage105[170]}
   );
   gpc1_1 gpc1_1_3412(
      {stage105[111]},
      {stage105[171]}
   );
   gpc1_1 gpc1_1_3413(
      {stage105[112]},
      {stage105[172]}
   );
   gpc1_1 gpc1_1_3414(
      {stage105[113]},
      {stage105[173]}
   );
   gpc1_1 gpc1_1_3415(
      {stage105[114]},
      {stage105[174]}
   );
   gpc1_1 gpc1_1_3416(
      {stage105[115]},
      {stage105[175]}
   );
   gpc1_1 gpc1_1_3417(
      {stage105[116]},
      {stage105[176]}
   );
   gpc1_1 gpc1_1_3418(
      {stage105[117]},
      {stage105[177]}
   );
   gpc1_1 gpc1_1_3419(
      {stage105[118]},
      {stage105[178]}
   );
   gpc1_1 gpc1_1_3420(
      {stage105[119]},
      {stage105[179]}
   );
   gpc1_1 gpc1_1_3421(
      {stage105[120]},
      {stage105[180]}
   );
   gpc1_1 gpc1_1_3422(
      {stage105[121]},
      {stage105[181]}
   );
   gpc606_5 gpc606_5_3423(
      {stage105[122], stage105[123], stage105[124], stage105[125], stage105[126], stage105[127]},
      {stage107[0], stage107[1], stage107[2], stage107[3], stage107[4], stage107[5]},
      {stage109[128], stage108[135], stage107[152], stage106[158], stage105[182]}
   );
   gpc1_1 gpc1_1_3424(
      {stage106[42]},
      {stage106[159]}
   );
   gpc1_1 gpc1_1_3425(
      {stage106[43]},
      {stage106[160]}
   );
   gpc1_1 gpc1_1_3426(
      {stage106[44]},
      {stage106[161]}
   );
   gpc1_1 gpc1_1_3427(
      {stage106[45]},
      {stage106[162]}
   );
   gpc1_1 gpc1_1_3428(
      {stage106[46]},
      {stage106[163]}
   );
   gpc1_1 gpc1_1_3429(
      {stage106[47]},
      {stage106[164]}
   );
   gpc1_1 gpc1_1_3430(
      {stage106[48]},
      {stage106[165]}
   );
   gpc1_1 gpc1_1_3431(
      {stage106[49]},
      {stage106[166]}
   );
   gpc1_1 gpc1_1_3432(
      {stage106[50]},
      {stage106[167]}
   );
   gpc1_1 gpc1_1_3433(
      {stage106[51]},
      {stage106[168]}
   );
   gpc1_1 gpc1_1_3434(
      {stage106[52]},
      {stage106[169]}
   );
   gpc1_1 gpc1_1_3435(
      {stage106[53]},
      {stage106[170]}
   );
   gpc1_1 gpc1_1_3436(
      {stage106[54]},
      {stage106[171]}
   );
   gpc1_1 gpc1_1_3437(
      {stage106[55]},
      {stage106[172]}
   );
   gpc1_1 gpc1_1_3438(
      {stage106[56]},
      {stage106[173]}
   );
   gpc1_1 gpc1_1_3439(
      {stage106[57]},
      {stage106[174]}
   );
   gpc1_1 gpc1_1_3440(
      {stage106[58]},
      {stage106[175]}
   );
   gpc1_1 gpc1_1_3441(
      {stage106[59]},
      {stage106[176]}
   );
   gpc1_1 gpc1_1_3442(
      {stage106[60]},
      {stage106[177]}
   );
   gpc1_1 gpc1_1_3443(
      {stage106[61]},
      {stage106[178]}
   );
   gpc1_1 gpc1_1_3444(
      {stage106[62]},
      {stage106[179]}
   );
   gpc1_1 gpc1_1_3445(
      {stage106[63]},
      {stage106[180]}
   );
   gpc1_1 gpc1_1_3446(
      {stage106[64]},
      {stage106[181]}
   );
   gpc1_1 gpc1_1_3447(
      {stage106[65]},
      {stage106[182]}
   );
   gpc1_1 gpc1_1_3448(
      {stage106[66]},
      {stage106[183]}
   );
   gpc1_1 gpc1_1_3449(
      {stage106[67]},
      {stage106[184]}
   );
   gpc615_5 gpc615_5_3450(
      {stage106[68], stage106[69], stage106[70], stage106[71], stage106[72]},
      {stage107[6]},
      {stage108[0], stage108[1], stage108[2], stage108[3], stage108[4], stage108[5]},
      {stage110[128], stage109[129], stage108[136], stage107[153], stage106[185]}
   );
   gpc615_5 gpc615_5_3451(
      {stage106[73], stage106[74], stage106[75], stage106[76], stage106[77]},
      {stage107[7]},
      {stage108[6], stage108[7], stage108[8], stage108[9], stage108[10], stage108[11]},
      {stage110[129], stage109[130], stage108[137], stage107[154], stage106[186]}
   );
   gpc615_5 gpc615_5_3452(
      {stage106[78], stage106[79], stage106[80], stage106[81], stage106[82]},
      {stage107[8]},
      {stage108[12], stage108[13], stage108[14], stage108[15], stage108[16], stage108[17]},
      {stage110[130], stage109[131], stage108[138], stage107[155], stage106[187]}
   );
   gpc615_5 gpc615_5_3453(
      {stage106[83], stage106[84], stage106[85], stage106[86], stage106[87]},
      {stage107[9]},
      {stage108[18], stage108[19], stage108[20], stage108[21], stage108[22], stage108[23]},
      {stage110[131], stage109[132], stage108[139], stage107[156], stage106[188]}
   );
   gpc615_5 gpc615_5_3454(
      {stage106[88], stage106[89], stage106[90], stage106[91], stage106[92]},
      {stage107[10]},
      {stage108[24], stage108[25], stage108[26], stage108[27], stage108[28], stage108[29]},
      {stage110[132], stage109[133], stage108[140], stage107[157], stage106[189]}
   );
   gpc615_5 gpc615_5_3455(
      {stage106[93], stage106[94], stage106[95], stage106[96], stage106[97]},
      {stage107[11]},
      {stage108[30], stage108[31], stage108[32], stage108[33], stage108[34], stage108[35]},
      {stage110[133], stage109[134], stage108[141], stage107[158], stage106[190]}
   );
   gpc615_5 gpc615_5_3456(
      {stage106[98], stage106[99], stage106[100], stage106[101], stage106[102]},
      {stage107[12]},
      {stage108[36], stage108[37], stage108[38], stage108[39], stage108[40], stage108[41]},
      {stage110[134], stage109[135], stage108[142], stage107[159], stage106[191]}
   );
   gpc615_5 gpc615_5_3457(
      {stage106[103], stage106[104], stage106[105], stage106[106], stage106[107]},
      {stage107[13]},
      {stage108[42], stage108[43], stage108[44], stage108[45], stage108[46], stage108[47]},
      {stage110[135], stage109[136], stage108[143], stage107[160], stage106[192]}
   );
   gpc615_5 gpc615_5_3458(
      {stage106[108], stage106[109], stage106[110], stage106[111], stage106[112]},
      {stage107[14]},
      {stage108[48], stage108[49], stage108[50], stage108[51], stage108[52], stage108[53]},
      {stage110[136], stage109[137], stage108[144], stage107[161], stage106[193]}
   );
   gpc615_5 gpc615_5_3459(
      {stage106[113], stage106[114], stage106[115], stage106[116], stage106[117]},
      {stage107[15]},
      {stage108[54], stage108[55], stage108[56], stage108[57], stage108[58], stage108[59]},
      {stage110[137], stage109[138], stage108[145], stage107[162], stage106[194]}
   );
   gpc615_5 gpc615_5_3460(
      {stage106[118], stage106[119], stage106[120], stage106[121], stage106[122]},
      {stage107[16]},
      {stage108[60], stage108[61], stage108[62], stage108[63], stage108[64], stage108[65]},
      {stage110[138], stage109[139], stage108[146], stage107[163], stage106[195]}
   );
   gpc615_5 gpc615_5_3461(
      {stage106[123], stage106[124], stage106[125], stage106[126], stage106[127]},
      {stage107[17]},
      {stage108[66], stage108[67], stage108[68], stage108[69], stage108[70], stage108[71]},
      {stage110[139], stage109[140], stage108[147], stage107[164], stage106[196]}
   );
   gpc1_1 gpc1_1_3462(
      {stage107[18]},
      {stage107[165]}
   );
   gpc1_1 gpc1_1_3463(
      {stage107[19]},
      {stage107[166]}
   );
   gpc1_1 gpc1_1_3464(
      {stage107[20]},
      {stage107[167]}
   );
   gpc1_1 gpc1_1_3465(
      {stage107[21]},
      {stage107[168]}
   );
   gpc606_5 gpc606_5_3466(
      {stage107[22], stage107[23], stage107[24], stage107[25], stage107[26], stage107[27]},
      {stage109[0], stage109[1], stage109[2], stage109[3], stage109[4], stage109[5]},
      {stage111[128], stage110[140], stage109[141], stage108[148], stage107[169]}
   );
   gpc606_5 gpc606_5_3467(
      {stage107[28], stage107[29], stage107[30], stage107[31], stage107[32], stage107[33]},
      {stage109[6], stage109[7], stage109[8], stage109[9], stage109[10], stage109[11]},
      {stage111[129], stage110[141], stage109[142], stage108[149], stage107[170]}
   );
   gpc606_5 gpc606_5_3468(
      {stage107[34], stage107[35], stage107[36], stage107[37], stage107[38], stage107[39]},
      {stage109[12], stage109[13], stage109[14], stage109[15], stage109[16], stage109[17]},
      {stage111[130], stage110[142], stage109[143], stage108[150], stage107[171]}
   );
   gpc606_5 gpc606_5_3469(
      {stage107[40], stage107[41], stage107[42], stage107[43], stage107[44], stage107[45]},
      {stage109[18], stage109[19], stage109[20], stage109[21], stage109[22], stage109[23]},
      {stage111[131], stage110[143], stage109[144], stage108[151], stage107[172]}
   );
   gpc606_5 gpc606_5_3470(
      {stage107[46], stage107[47], stage107[48], stage107[49], stage107[50], stage107[51]},
      {stage109[24], stage109[25], stage109[26], stage109[27], stage109[28], stage109[29]},
      {stage111[132], stage110[144], stage109[145], stage108[152], stage107[173]}
   );
   gpc606_5 gpc606_5_3471(
      {stage107[52], stage107[53], stage107[54], stage107[55], stage107[56], stage107[57]},
      {stage109[30], stage109[31], stage109[32], stage109[33], stage109[34], stage109[35]},
      {stage111[133], stage110[145], stage109[146], stage108[153], stage107[174]}
   );
   gpc606_5 gpc606_5_3472(
      {stage107[58], stage107[59], stage107[60], stage107[61], stage107[62], stage107[63]},
      {stage109[36], stage109[37], stage109[38], stage109[39], stage109[40], stage109[41]},
      {stage111[134], stage110[146], stage109[147], stage108[154], stage107[175]}
   );
   gpc606_5 gpc606_5_3473(
      {stage107[64], stage107[65], stage107[66], stage107[67], stage107[68], stage107[69]},
      {stage109[42], stage109[43], stage109[44], stage109[45], stage109[46], stage109[47]},
      {stage111[135], stage110[147], stage109[148], stage108[155], stage107[176]}
   );
   gpc606_5 gpc606_5_3474(
      {stage107[70], stage107[71], stage107[72], stage107[73], stage107[74], stage107[75]},
      {stage109[48], stage109[49], stage109[50], stage109[51], stage109[52], stage109[53]},
      {stage111[136], stage110[148], stage109[149], stage108[156], stage107[177]}
   );
   gpc606_5 gpc606_5_3475(
      {stage107[76], stage107[77], stage107[78], stage107[79], stage107[80], stage107[81]},
      {stage109[54], stage109[55], stage109[56], stage109[57], stage109[58], stage109[59]},
      {stage111[137], stage110[149], stage109[150], stage108[157], stage107[178]}
   );
   gpc606_5 gpc606_5_3476(
      {stage107[82], stage107[83], stage107[84], stage107[85], stage107[86], stage107[87]},
      {stage109[60], stage109[61], stage109[62], stage109[63], stage109[64], stage109[65]},
      {stage111[138], stage110[150], stage109[151], stage108[158], stage107[179]}
   );
   gpc606_5 gpc606_5_3477(
      {stage107[88], stage107[89], stage107[90], stage107[91], stage107[92], stage107[93]},
      {stage109[66], stage109[67], stage109[68], stage109[69], stage109[70], stage109[71]},
      {stage111[139], stage110[151], stage109[152], stage108[159], stage107[180]}
   );
   gpc606_5 gpc606_5_3478(
      {stage107[94], stage107[95], stage107[96], stage107[97], stage107[98], stage107[99]},
      {stage109[72], stage109[73], stage109[74], stage109[75], stage109[76], stage109[77]},
      {stage111[140], stage110[152], stage109[153], stage108[160], stage107[181]}
   );
   gpc606_5 gpc606_5_3479(
      {stage107[100], stage107[101], stage107[102], stage107[103], stage107[104], stage107[105]},
      {stage109[78], stage109[79], stage109[80], stage109[81], stage109[82], stage109[83]},
      {stage111[141], stage110[153], stage109[154], stage108[161], stage107[182]}
   );
   gpc606_5 gpc606_5_3480(
      {stage107[106], stage107[107], stage107[108], stage107[109], stage107[110], stage107[111]},
      {stage109[84], stage109[85], stage109[86], stage109[87], stage109[88], stage109[89]},
      {stage111[142], stage110[154], stage109[155], stage108[162], stage107[183]}
   );
   gpc606_5 gpc606_5_3481(
      {stage107[112], stage107[113], stage107[114], stage107[115], stage107[116], stage107[117]},
      {stage109[90], stage109[91], stage109[92], stage109[93], stage109[94], stage109[95]},
      {stage111[143], stage110[155], stage109[156], stage108[163], stage107[184]}
   );
   gpc615_5 gpc615_5_3482(
      {stage107[118], stage107[119], stage107[120], stage107[121], stage107[122]},
      {stage108[72]},
      {stage109[96], stage109[97], stage109[98], stage109[99], stage109[100], stage109[101]},
      {stage111[144], stage110[156], stage109[157], stage108[164], stage107[185]}
   );
   gpc615_5 gpc615_5_3483(
      {stage107[123], stage107[124], stage107[125], stage107[126], stage107[127]},
      {stage108[73]},
      {stage109[102], stage109[103], stage109[104], stage109[105], stage109[106], stage109[107]},
      {stage111[145], stage110[157], stage109[158], stage108[165], stage107[186]}
   );
   gpc1_1 gpc1_1_3484(
      {stage108[74]},
      {stage108[166]}
   );
   gpc1_1 gpc1_1_3485(
      {stage108[75]},
      {stage108[167]}
   );
   gpc1_1 gpc1_1_3486(
      {stage108[76]},
      {stage108[168]}
   );
   gpc1_1 gpc1_1_3487(
      {stage108[77]},
      {stage108[169]}
   );
   gpc1_1 gpc1_1_3488(
      {stage108[78]},
      {stage108[170]}
   );
   gpc1_1 gpc1_1_3489(
      {stage108[79]},
      {stage108[171]}
   );
   gpc606_5 gpc606_5_3490(
      {stage108[80], stage108[81], stage108[82], stage108[83], stage108[84], stage108[85]},
      {stage110[0], stage110[1], stage110[2], stage110[3], stage110[4], stage110[5]},
      {stage112[128], stage111[146], stage110[158], stage109[159], stage108[172]}
   );
   gpc606_5 gpc606_5_3491(
      {stage108[86], stage108[87], stage108[88], stage108[89], stage108[90], stage108[91]},
      {stage110[6], stage110[7], stage110[8], stage110[9], stage110[10], stage110[11]},
      {stage112[129], stage111[147], stage110[159], stage109[160], stage108[173]}
   );
   gpc606_5 gpc606_5_3492(
      {stage108[92], stage108[93], stage108[94], stage108[95], stage108[96], stage108[97]},
      {stage110[12], stage110[13], stage110[14], stage110[15], stage110[16], stage110[17]},
      {stage112[130], stage111[148], stage110[160], stage109[161], stage108[174]}
   );
   gpc606_5 gpc606_5_3493(
      {stage108[98], stage108[99], stage108[100], stage108[101], stage108[102], stage108[103]},
      {stage110[18], stage110[19], stage110[20], stage110[21], stage110[22], stage110[23]},
      {stage112[131], stage111[149], stage110[161], stage109[162], stage108[175]}
   );
   gpc606_5 gpc606_5_3494(
      {stage108[104], stage108[105], stage108[106], stage108[107], stage108[108], stage108[109]},
      {stage110[24], stage110[25], stage110[26], stage110[27], stage110[28], stage110[29]},
      {stage112[132], stage111[150], stage110[162], stage109[163], stage108[176]}
   );
   gpc606_5 gpc606_5_3495(
      {stage108[110], stage108[111], stage108[112], stage108[113], stage108[114], stage108[115]},
      {stage110[30], stage110[31], stage110[32], stage110[33], stage110[34], stage110[35]},
      {stage112[133], stage111[151], stage110[163], stage109[164], stage108[177]}
   );
   gpc606_5 gpc606_5_3496(
      {stage108[116], stage108[117], stage108[118], stage108[119], stage108[120], stage108[121]},
      {stage110[36], stage110[37], stage110[38], stage110[39], stage110[40], stage110[41]},
      {stage112[134], stage111[152], stage110[164], stage109[165], stage108[178]}
   );
   gpc606_5 gpc606_5_3497(
      {stage108[122], stage108[123], stage108[124], stage108[125], stage108[126], stage108[127]},
      {stage110[42], stage110[43], stage110[44], stage110[45], stage110[46], stage110[47]},
      {stage112[135], stage111[153], stage110[165], stage109[166], stage108[179]}
   );
   gpc1_1 gpc1_1_3498(
      {stage109[108]},
      {stage109[167]}
   );
   gpc1_1 gpc1_1_3499(
      {stage109[109]},
      {stage109[168]}
   );
   gpc1_1 gpc1_1_3500(
      {stage109[110]},
      {stage109[169]}
   );
   gpc1_1 gpc1_1_3501(
      {stage109[111]},
      {stage109[170]}
   );
   gpc1_1 gpc1_1_3502(
      {stage109[112]},
      {stage109[171]}
   );
   gpc1_1 gpc1_1_3503(
      {stage109[113]},
      {stage109[172]}
   );
   gpc1_1 gpc1_1_3504(
      {stage109[114]},
      {stage109[173]}
   );
   gpc1_1 gpc1_1_3505(
      {stage109[115]},
      {stage109[174]}
   );
   gpc1_1 gpc1_1_3506(
      {stage109[116]},
      {stage109[175]}
   );
   gpc1_1 gpc1_1_3507(
      {stage109[117]},
      {stage109[176]}
   );
   gpc1_1 gpc1_1_3508(
      {stage109[118]},
      {stage109[177]}
   );
   gpc1_1 gpc1_1_3509(
      {stage109[119]},
      {stage109[178]}
   );
   gpc1_1 gpc1_1_3510(
      {stage109[120]},
      {stage109[179]}
   );
   gpc1_1 gpc1_1_3511(
      {stage109[121]},
      {stage109[180]}
   );
   gpc1_1 gpc1_1_3512(
      {stage109[122]},
      {stage109[181]}
   );
   gpc615_5 gpc615_5_3513(
      {stage109[123], stage109[124], stage109[125], stage109[126], stage109[127]},
      {stage110[48]},
      {stage111[0], stage111[1], stage111[2], stage111[3], stage111[4], stage111[5]},
      {stage113[128], stage112[136], stage111[154], stage110[166], stage109[182]}
   );
   gpc1_1 gpc1_1_3514(
      {stage110[49]},
      {stage110[167]}
   );
   gpc1_1 gpc1_1_3515(
      {stage110[50]},
      {stage110[168]}
   );
   gpc1_1 gpc1_1_3516(
      {stage110[51]},
      {stage110[169]}
   );
   gpc1_1 gpc1_1_3517(
      {stage110[52]},
      {stage110[170]}
   );
   gpc1_1 gpc1_1_3518(
      {stage110[53]},
      {stage110[171]}
   );
   gpc1_1 gpc1_1_3519(
      {stage110[54]},
      {stage110[172]}
   );
   gpc1_1 gpc1_1_3520(
      {stage110[55]},
      {stage110[173]}
   );
   gpc1_1 gpc1_1_3521(
      {stage110[56]},
      {stage110[174]}
   );
   gpc1_1 gpc1_1_3522(
      {stage110[57]},
      {stage110[175]}
   );
   gpc1_1 gpc1_1_3523(
      {stage110[58]},
      {stage110[176]}
   );
   gpc1_1 gpc1_1_3524(
      {stage110[59]},
      {stage110[177]}
   );
   gpc1_1 gpc1_1_3525(
      {stage110[60]},
      {stage110[178]}
   );
   gpc1_1 gpc1_1_3526(
      {stage110[61]},
      {stage110[179]}
   );
   gpc1_1 gpc1_1_3527(
      {stage110[62]},
      {stage110[180]}
   );
   gpc1_1 gpc1_1_3528(
      {stage110[63]},
      {stage110[181]}
   );
   gpc1_1 gpc1_1_3529(
      {stage110[64]},
      {stage110[182]}
   );
   gpc1_1 gpc1_1_3530(
      {stage110[65]},
      {stage110[183]}
   );
   gpc1_1 gpc1_1_3531(
      {stage110[66]},
      {stage110[184]}
   );
   gpc1_1 gpc1_1_3532(
      {stage110[67]},
      {stage110[185]}
   );
   gpc1_1 gpc1_1_3533(
      {stage110[68]},
      {stage110[186]}
   );
   gpc1_1 gpc1_1_3534(
      {stage110[69]},
      {stage110[187]}
   );
   gpc606_5 gpc606_5_3535(
      {stage110[70], stage110[71], stage110[72], stage110[73], stage110[74], stage110[75]},
      {stage112[0], stage112[1], stage112[2], stage112[3], stage112[4], stage112[5]},
      {stage114[128], stage113[129], stage112[137], stage111[155], stage110[188]}
   );
   gpc606_5 gpc606_5_3536(
      {stage110[76], stage110[77], stage110[78], stage110[79], stage110[80], stage110[81]},
      {stage112[6], stage112[7], stage112[8], stage112[9], stage112[10], stage112[11]},
      {stage114[129], stage113[130], stage112[138], stage111[156], stage110[189]}
   );
   gpc606_5 gpc606_5_3537(
      {stage110[82], stage110[83], stage110[84], stage110[85], stage110[86], stage110[87]},
      {stage112[12], stage112[13], stage112[14], stage112[15], stage112[16], stage112[17]},
      {stage114[130], stage113[131], stage112[139], stage111[157], stage110[190]}
   );
   gpc615_5 gpc615_5_3538(
      {stage110[88], stage110[89], stage110[90], stage110[91], stage110[92]},
      {stage111[6]},
      {stage112[18], stage112[19], stage112[20], stage112[21], stage112[22], stage112[23]},
      {stage114[131], stage113[132], stage112[140], stage111[158], stage110[191]}
   );
   gpc615_5 gpc615_5_3539(
      {stage110[93], stage110[94], stage110[95], stage110[96], stage110[97]},
      {stage111[7]},
      {stage112[24], stage112[25], stage112[26], stage112[27], stage112[28], stage112[29]},
      {stage114[132], stage113[133], stage112[141], stage111[159], stage110[192]}
   );
   gpc615_5 gpc615_5_3540(
      {stage110[98], stage110[99], stage110[100], stage110[101], stage110[102]},
      {stage111[8]},
      {stage112[30], stage112[31], stage112[32], stage112[33], stage112[34], stage112[35]},
      {stage114[133], stage113[134], stage112[142], stage111[160], stage110[193]}
   );
   gpc615_5 gpc615_5_3541(
      {stage110[103], stage110[104], stage110[105], stage110[106], stage110[107]},
      {stage111[9]},
      {stage112[36], stage112[37], stage112[38], stage112[39], stage112[40], stage112[41]},
      {stage114[134], stage113[135], stage112[143], stage111[161], stage110[194]}
   );
   gpc615_5 gpc615_5_3542(
      {stage110[108], stage110[109], stage110[110], stage110[111], stage110[112]},
      {stage111[10]},
      {stage112[42], stage112[43], stage112[44], stage112[45], stage112[46], stage112[47]},
      {stage114[135], stage113[136], stage112[144], stage111[162], stage110[195]}
   );
   gpc615_5 gpc615_5_3543(
      {stage110[113], stage110[114], stage110[115], stage110[116], stage110[117]},
      {stage111[11]},
      {stage112[48], stage112[49], stage112[50], stage112[51], stage112[52], stage112[53]},
      {stage114[136], stage113[137], stage112[145], stage111[163], stage110[196]}
   );
   gpc615_5 gpc615_5_3544(
      {stage110[118], stage110[119], stage110[120], stage110[121], stage110[122]},
      {stage111[12]},
      {stage112[54], stage112[55], stage112[56], stage112[57], stage112[58], stage112[59]},
      {stage114[137], stage113[138], stage112[146], stage111[164], stage110[197]}
   );
   gpc615_5 gpc615_5_3545(
      {stage110[123], stage110[124], stage110[125], stage110[126], stage110[127]},
      {stage111[13]},
      {stage112[60], stage112[61], stage112[62], stage112[63], stage112[64], stage112[65]},
      {stage114[138], stage113[139], stage112[147], stage111[165], stage110[198]}
   );
   gpc1_1 gpc1_1_3546(
      {stage111[14]},
      {stage111[166]}
   );
   gpc1_1 gpc1_1_3547(
      {stage111[15]},
      {stage111[167]}
   );
   gpc1_1 gpc1_1_3548(
      {stage111[16]},
      {stage111[168]}
   );
   gpc1_1 gpc1_1_3549(
      {stage111[17]},
      {stage111[169]}
   );
   gpc1_1 gpc1_1_3550(
      {stage111[18]},
      {stage111[170]}
   );
   gpc1_1 gpc1_1_3551(
      {stage111[19]},
      {stage111[171]}
   );
   gpc1_1 gpc1_1_3552(
      {stage111[20]},
      {stage111[172]}
   );
   gpc1_1 gpc1_1_3553(
      {stage111[21]},
      {stage111[173]}
   );
   gpc1_1 gpc1_1_3554(
      {stage111[22]},
      {stage111[174]}
   );
   gpc1_1 gpc1_1_3555(
      {stage111[23]},
      {stage111[175]}
   );
   gpc1_1 gpc1_1_3556(
      {stage111[24]},
      {stage111[176]}
   );
   gpc1_1 gpc1_1_3557(
      {stage111[25]},
      {stage111[177]}
   );
   gpc1_1 gpc1_1_3558(
      {stage111[26]},
      {stage111[178]}
   );
   gpc1_1 gpc1_1_3559(
      {stage111[27]},
      {stage111[179]}
   );
   gpc1_1 gpc1_1_3560(
      {stage111[28]},
      {stage111[180]}
   );
   gpc1_1 gpc1_1_3561(
      {stage111[29]},
      {stage111[181]}
   );
   gpc1_1 gpc1_1_3562(
      {stage111[30]},
      {stage111[182]}
   );
   gpc1_1 gpc1_1_3563(
      {stage111[31]},
      {stage111[183]}
   );
   gpc1_1 gpc1_1_3564(
      {stage111[32]},
      {stage111[184]}
   );
   gpc1_1 gpc1_1_3565(
      {stage111[33]},
      {stage111[185]}
   );
   gpc1_1 gpc1_1_3566(
      {stage111[34]},
      {stage111[186]}
   );
   gpc1_1 gpc1_1_3567(
      {stage111[35]},
      {stage111[187]}
   );
   gpc1_1 gpc1_1_3568(
      {stage111[36]},
      {stage111[188]}
   );
   gpc1_1 gpc1_1_3569(
      {stage111[37]},
      {stage111[189]}
   );
   gpc1_1 gpc1_1_3570(
      {stage111[38]},
      {stage111[190]}
   );
   gpc1_1 gpc1_1_3571(
      {stage111[39]},
      {stage111[191]}
   );
   gpc1_1 gpc1_1_3572(
      {stage111[40]},
      {stage111[192]}
   );
   gpc1_1 gpc1_1_3573(
      {stage111[41]},
      {stage111[193]}
   );
   gpc1_1 gpc1_1_3574(
      {stage111[42]},
      {stage111[194]}
   );
   gpc1_1 gpc1_1_3575(
      {stage111[43]},
      {stage111[195]}
   );
   gpc1_1 gpc1_1_3576(
      {stage111[44]},
      {stage111[196]}
   );
   gpc1_1 gpc1_1_3577(
      {stage111[45]},
      {stage111[197]}
   );
   gpc1_1 gpc1_1_3578(
      {stage111[46]},
      {stage111[198]}
   );
   gpc1_1 gpc1_1_3579(
      {stage111[47]},
      {stage111[199]}
   );
   gpc1_1 gpc1_1_3580(
      {stage111[48]},
      {stage111[200]}
   );
   gpc1_1 gpc1_1_3581(
      {stage111[49]},
      {stage111[201]}
   );
   gpc606_5 gpc606_5_3582(
      {stage111[50], stage111[51], stage111[52], stage111[53], stage111[54], stage111[55]},
      {stage113[0], stage113[1], stage113[2], stage113[3], stage113[4], stage113[5]},
      {stage115[128], stage114[139], stage113[140], stage112[148], stage111[202]}
   );
   gpc606_5 gpc606_5_3583(
      {stage111[56], stage111[57], stage111[58], stage111[59], stage111[60], stage111[61]},
      {stage113[6], stage113[7], stage113[8], stage113[9], stage113[10], stage113[11]},
      {stage115[129], stage114[140], stage113[141], stage112[149], stage111[203]}
   );
   gpc606_5 gpc606_5_3584(
      {stage111[62], stage111[63], stage111[64], stage111[65], stage111[66], stage111[67]},
      {stage113[12], stage113[13], stage113[14], stage113[15], stage113[16], stage113[17]},
      {stage115[130], stage114[141], stage113[142], stage112[150], stage111[204]}
   );
   gpc606_5 gpc606_5_3585(
      {stage111[68], stage111[69], stage111[70], stage111[71], stage111[72], stage111[73]},
      {stage113[18], stage113[19], stage113[20], stage113[21], stage113[22], stage113[23]},
      {stage115[131], stage114[142], stage113[143], stage112[151], stage111[205]}
   );
   gpc606_5 gpc606_5_3586(
      {stage111[74], stage111[75], stage111[76], stage111[77], stage111[78], stage111[79]},
      {stage113[24], stage113[25], stage113[26], stage113[27], stage113[28], stage113[29]},
      {stage115[132], stage114[143], stage113[144], stage112[152], stage111[206]}
   );
   gpc606_5 gpc606_5_3587(
      {stage111[80], stage111[81], stage111[82], stage111[83], stage111[84], stage111[85]},
      {stage113[30], stage113[31], stage113[32], stage113[33], stage113[34], stage113[35]},
      {stage115[133], stage114[144], stage113[145], stage112[153], stage111[207]}
   );
   gpc606_5 gpc606_5_3588(
      {stage111[86], stage111[87], stage111[88], stage111[89], stage111[90], stage111[91]},
      {stage113[36], stage113[37], stage113[38], stage113[39], stage113[40], stage113[41]},
      {stage115[134], stage114[145], stage113[146], stage112[154], stage111[208]}
   );
   gpc606_5 gpc606_5_3589(
      {stage111[92], stage111[93], stage111[94], stage111[95], stage111[96], stage111[97]},
      {stage113[42], stage113[43], stage113[44], stage113[45], stage113[46], stage113[47]},
      {stage115[135], stage114[146], stage113[147], stage112[155], stage111[209]}
   );
   gpc606_5 gpc606_5_3590(
      {stage111[98], stage111[99], stage111[100], stage111[101], stage111[102], stage111[103]},
      {stage113[48], stage113[49], stage113[50], stage113[51], stage113[52], stage113[53]},
      {stage115[136], stage114[147], stage113[148], stage112[156], stage111[210]}
   );
   gpc606_5 gpc606_5_3591(
      {stage111[104], stage111[105], stage111[106], stage111[107], stage111[108], stage111[109]},
      {stage113[54], stage113[55], stage113[56], stage113[57], stage113[58], stage113[59]},
      {stage115[137], stage114[148], stage113[149], stage112[157], stage111[211]}
   );
   gpc606_5 gpc606_5_3592(
      {stage111[110], stage111[111], stage111[112], stage111[113], stage111[114], stage111[115]},
      {stage113[60], stage113[61], stage113[62], stage113[63], stage113[64], stage113[65]},
      {stage115[138], stage114[149], stage113[150], stage112[158], stage111[212]}
   );
   gpc606_5 gpc606_5_3593(
      {stage111[116], stage111[117], stage111[118], stage111[119], stage111[120], stage111[121]},
      {stage113[66], stage113[67], stage113[68], stage113[69], stage113[70], stage113[71]},
      {stage115[139], stage114[150], stage113[151], stage112[159], stage111[213]}
   );
   gpc606_5 gpc606_5_3594(
      {stage111[122], stage111[123], stage111[124], stage111[125], stage111[126], stage111[127]},
      {stage113[72], stage113[73], stage113[74], stage113[75], stage113[76], stage113[77]},
      {stage115[140], stage114[151], stage113[152], stage112[160], stage111[214]}
   );
   gpc1_1 gpc1_1_3595(
      {stage112[66]},
      {stage112[161]}
   );
   gpc1_1 gpc1_1_3596(
      {stage112[67]},
      {stage112[162]}
   );
   gpc1_1 gpc1_1_3597(
      {stage112[68]},
      {stage112[163]}
   );
   gpc1_1 gpc1_1_3598(
      {stage112[69]},
      {stage112[164]}
   );
   gpc1_1 gpc1_1_3599(
      {stage112[70]},
      {stage112[165]}
   );
   gpc1_1 gpc1_1_3600(
      {stage112[71]},
      {stage112[166]}
   );
   gpc1_1 gpc1_1_3601(
      {stage112[72]},
      {stage112[167]}
   );
   gpc1_1 gpc1_1_3602(
      {stage112[73]},
      {stage112[168]}
   );
   gpc1_1 gpc1_1_3603(
      {stage112[74]},
      {stage112[169]}
   );
   gpc1_1 gpc1_1_3604(
      {stage112[75]},
      {stage112[170]}
   );
   gpc1_1 gpc1_1_3605(
      {stage112[76]},
      {stage112[171]}
   );
   gpc1_1 gpc1_1_3606(
      {stage112[77]},
      {stage112[172]}
   );
   gpc1_1 gpc1_1_3607(
      {stage112[78]},
      {stage112[173]}
   );
   gpc1_1 gpc1_1_3608(
      {stage112[79]},
      {stage112[174]}
   );
   gpc1_1 gpc1_1_3609(
      {stage112[80]},
      {stage112[175]}
   );
   gpc1_1 gpc1_1_3610(
      {stage112[81]},
      {stage112[176]}
   );
   gpc1_1 gpc1_1_3611(
      {stage112[82]},
      {stage112[177]}
   );
   gpc1_1 gpc1_1_3612(
      {stage112[83]},
      {stage112[178]}
   );
   gpc1_1 gpc1_1_3613(
      {stage112[84]},
      {stage112[179]}
   );
   gpc1_1 gpc1_1_3614(
      {stage112[85]},
      {stage112[180]}
   );
   gpc1_1 gpc1_1_3615(
      {stage112[86]},
      {stage112[181]}
   );
   gpc1_1 gpc1_1_3616(
      {stage112[87]},
      {stage112[182]}
   );
   gpc1_1 gpc1_1_3617(
      {stage112[88]},
      {stage112[183]}
   );
   gpc1_1 gpc1_1_3618(
      {stage112[89]},
      {stage112[184]}
   );
   gpc606_5 gpc606_5_3619(
      {stage112[90], stage112[91], stage112[92], stage112[93], stage112[94], stage112[95]},
      {stage114[0], stage114[1], stage114[2], stage114[3], stage114[4], stage114[5]},
      {stage116[128], stage115[141], stage114[152], stage113[153], stage112[185]}
   );
   gpc606_5 gpc606_5_3620(
      {stage112[96], stage112[97], stage112[98], stage112[99], stage112[100], stage112[101]},
      {stage114[6], stage114[7], stage114[8], stage114[9], stage114[10], stage114[11]},
      {stage116[129], stage115[142], stage114[153], stage113[154], stage112[186]}
   );
   gpc606_5 gpc606_5_3621(
      {stage112[102], stage112[103], stage112[104], stage112[105], stage112[106], stage112[107]},
      {stage114[12], stage114[13], stage114[14], stage114[15], stage114[16], stage114[17]},
      {stage116[130], stage115[143], stage114[154], stage113[155], stage112[187]}
   );
   gpc606_5 gpc606_5_3622(
      {stage112[108], stage112[109], stage112[110], stage112[111], stage112[112], stage112[113]},
      {stage114[18], stage114[19], stage114[20], stage114[21], stage114[22], stage114[23]},
      {stage116[131], stage115[144], stage114[155], stage113[156], stage112[188]}
   );
   gpc606_5 gpc606_5_3623(
      {stage112[114], stage112[115], stage112[116], stage112[117], stage112[118], stage112[119]},
      {stage114[24], stage114[25], stage114[26], stage114[27], stage114[28], stage114[29]},
      {stage116[132], stage115[145], stage114[156], stage113[157], stage112[189]}
   );
   gpc1343_5 gpc1343_5_3624(
      {stage112[120], stage112[121], stage112[122]},
      {stage113[78], stage113[79], stage113[80], stage113[81]},
      {stage114[30], stage114[31], stage114[32]},
      {stage115[0]},
      {stage116[133], stage115[146], stage114[157], stage113[158], stage112[190]}
   );
   gpc2135_5 gpc2135_5_3625(
      {stage112[123], stage112[124], stage112[125], stage112[126], stage112[127]},
      {stage113[82], stage113[83], stage113[84]},
      {stage114[33]},
      {stage115[1], stage115[2]},
      {stage116[134], stage115[147], stage114[158], stage113[159], stage112[191]}
   );
   gpc1_1 gpc1_1_3626(
      {stage113[85]},
      {stage113[160]}
   );
   gpc1_1 gpc1_1_3627(
      {stage113[86]},
      {stage113[161]}
   );
   gpc1_1 gpc1_1_3628(
      {stage113[87]},
      {stage113[162]}
   );
   gpc1_1 gpc1_1_3629(
      {stage113[88]},
      {stage113[163]}
   );
   gpc1_1 gpc1_1_3630(
      {stage113[89]},
      {stage113[164]}
   );
   gpc1_1 gpc1_1_3631(
      {stage113[90]},
      {stage113[165]}
   );
   gpc1_1 gpc1_1_3632(
      {stage113[91]},
      {stage113[166]}
   );
   gpc1_1 gpc1_1_3633(
      {stage113[92]},
      {stage113[167]}
   );
   gpc1_1 gpc1_1_3634(
      {stage113[93]},
      {stage113[168]}
   );
   gpc1_1 gpc1_1_3635(
      {stage113[94]},
      {stage113[169]}
   );
   gpc1_1 gpc1_1_3636(
      {stage113[95]},
      {stage113[170]}
   );
   gpc1_1 gpc1_1_3637(
      {stage113[96]},
      {stage113[171]}
   );
   gpc1_1 gpc1_1_3638(
      {stage113[97]},
      {stage113[172]}
   );
   gpc1_1 gpc1_1_3639(
      {stage113[98]},
      {stage113[173]}
   );
   gpc1_1 gpc1_1_3640(
      {stage113[99]},
      {stage113[174]}
   );
   gpc1_1 gpc1_1_3641(
      {stage113[100]},
      {stage113[175]}
   );
   gpc1_1 gpc1_1_3642(
      {stage113[101]},
      {stage113[176]}
   );
   gpc1_1 gpc1_1_3643(
      {stage113[102]},
      {stage113[177]}
   );
   gpc1_1 gpc1_1_3644(
      {stage113[103]},
      {stage113[178]}
   );
   gpc606_5 gpc606_5_3645(
      {stage113[104], stage113[105], stage113[106], stage113[107], stage113[108], stage113[109]},
      {stage115[3], stage115[4], stage115[5], stage115[6], stage115[7], stage115[8]},
      {stage117[128], stage116[135], stage115[148], stage114[159], stage113[179]}
   );
   gpc606_5 gpc606_5_3646(
      {stage113[110], stage113[111], stage113[112], stage113[113], stage113[114], stage113[115]},
      {stage115[9], stage115[10], stage115[11], stage115[12], stage115[13], stage115[14]},
      {stage117[129], stage116[136], stage115[149], stage114[160], stage113[180]}
   );
   gpc606_5 gpc606_5_3647(
      {stage113[116], stage113[117], stage113[118], stage113[119], stage113[120], stage113[121]},
      {stage115[15], stage115[16], stage115[17], stage115[18], stage115[19], stage115[20]},
      {stage117[130], stage116[137], stage115[150], stage114[161], stage113[181]}
   );
   gpc606_5 gpc606_5_3648(
      {stage113[122], stage113[123], stage113[124], stage113[125], stage113[126], stage113[127]},
      {stage115[21], stage115[22], stage115[23], stage115[24], stage115[25], stage115[26]},
      {stage117[131], stage116[138], stage115[151], stage114[162], stage113[182]}
   );
   gpc1_1 gpc1_1_3649(
      {stage114[34]},
      {stage114[163]}
   );
   gpc1_1 gpc1_1_3650(
      {stage114[35]},
      {stage114[164]}
   );
   gpc1_1 gpc1_1_3651(
      {stage114[36]},
      {stage114[165]}
   );
   gpc1_1 gpc1_1_3652(
      {stage114[37]},
      {stage114[166]}
   );
   gpc1_1 gpc1_1_3653(
      {stage114[38]},
      {stage114[167]}
   );
   gpc1_1 gpc1_1_3654(
      {stage114[39]},
      {stage114[168]}
   );
   gpc1_1 gpc1_1_3655(
      {stage114[40]},
      {stage114[169]}
   );
   gpc606_5 gpc606_5_3656(
      {stage114[41], stage114[42], stage114[43], stage114[44], stage114[45], stage114[46]},
      {stage116[0], stage116[1], stage116[2], stage116[3], stage116[4], stage116[5]},
      {stage118[128], stage117[132], stage116[139], stage115[152], stage114[170]}
   );
   gpc606_5 gpc606_5_3657(
      {stage114[47], stage114[48], stage114[49], stage114[50], stage114[51], stage114[52]},
      {stage116[6], stage116[7], stage116[8], stage116[9], stage116[10], stage116[11]},
      {stage118[129], stage117[133], stage116[140], stage115[153], stage114[171]}
   );
   gpc606_5 gpc606_5_3658(
      {stage114[53], stage114[54], stage114[55], stage114[56], stage114[57], stage114[58]},
      {stage116[12], stage116[13], stage116[14], stage116[15], stage116[16], stage116[17]},
      {stage118[130], stage117[134], stage116[141], stage115[154], stage114[172]}
   );
   gpc606_5 gpc606_5_3659(
      {stage114[59], stage114[60], stage114[61], stage114[62], stage114[63], stage114[64]},
      {stage116[18], stage116[19], stage116[20], stage116[21], stage116[22], stage116[23]},
      {stage118[131], stage117[135], stage116[142], stage115[155], stage114[173]}
   );
   gpc207_4 gpc207_4_3660(
      {stage114[65], stage114[66], stage114[67], stage114[68], stage114[69], stage114[70], stage114[71]},
      {stage116[24], stage116[25]},
      {stage117[136], stage116[143], stage115[156], stage114[174]}
   );
   gpc207_4 gpc207_4_3661(
      {stage114[72], stage114[73], stage114[74], stage114[75], stage114[76], stage114[77], stage114[78]},
      {stage116[26], stage116[27]},
      {stage117[137], stage116[144], stage115[157], stage114[175]}
   );
   gpc207_4 gpc207_4_3662(
      {stage114[79], stage114[80], stage114[81], stage114[82], stage114[83], stage114[84], stage114[85]},
      {stage116[28], stage116[29]},
      {stage117[138], stage116[145], stage115[158], stage114[176]}
   );
   gpc207_4 gpc207_4_3663(
      {stage114[86], stage114[87], stage114[88], stage114[89], stage114[90], stage114[91], stage114[92]},
      {stage116[30], stage116[31]},
      {stage117[139], stage116[146], stage115[159], stage114[177]}
   );
   gpc207_4 gpc207_4_3664(
      {stage114[93], stage114[94], stage114[95], stage114[96], stage114[97], stage114[98], stage114[99]},
      {stage116[32], stage116[33]},
      {stage117[140], stage116[147], stage115[160], stage114[178]}
   );
   gpc207_4 gpc207_4_3665(
      {stage114[100], stage114[101], stage114[102], stage114[103], stage114[104], stage114[105], stage114[106]},
      {stage116[34], stage116[35]},
      {stage117[141], stage116[148], stage115[161], stage114[179]}
   );
   gpc207_4 gpc207_4_3666(
      {stage114[107], stage114[108], stage114[109], stage114[110], stage114[111], stage114[112], stage114[113]},
      {stage116[36], stage116[37]},
      {stage117[142], stage116[149], stage115[162], stage114[180]}
   );
   gpc207_4 gpc207_4_3667(
      {stage114[114], stage114[115], stage114[116], stage114[117], stage114[118], stage114[119], stage114[120]},
      {stage116[38], stage116[39]},
      {stage117[143], stage116[150], stage115[163], stage114[181]}
   );
   gpc207_4 gpc207_4_3668(
      {stage114[121], stage114[122], stage114[123], stage114[124], stage114[125], stage114[126], stage114[127]},
      {stage116[40], stage116[41]},
      {stage117[144], stage116[151], stage115[164], stage114[182]}
   );
   gpc1_1 gpc1_1_3669(
      {stage115[27]},
      {stage115[165]}
   );
   gpc1_1 gpc1_1_3670(
      {stage115[28]},
      {stage115[166]}
   );
   gpc1_1 gpc1_1_3671(
      {stage115[29]},
      {stage115[167]}
   );
   gpc1_1 gpc1_1_3672(
      {stage115[30]},
      {stage115[168]}
   );
   gpc1_1 gpc1_1_3673(
      {stage115[31]},
      {stage115[169]}
   );
   gpc1_1 gpc1_1_3674(
      {stage115[32]},
      {stage115[170]}
   );
   gpc1_1 gpc1_1_3675(
      {stage115[33]},
      {stage115[171]}
   );
   gpc1_1 gpc1_1_3676(
      {stage115[34]},
      {stage115[172]}
   );
   gpc1_1 gpc1_1_3677(
      {stage115[35]},
      {stage115[173]}
   );
   gpc1_1 gpc1_1_3678(
      {stage115[36]},
      {stage115[174]}
   );
   gpc1_1 gpc1_1_3679(
      {stage115[37]},
      {stage115[175]}
   );
   gpc1_1 gpc1_1_3680(
      {stage115[38]},
      {stage115[176]}
   );
   gpc1_1 gpc1_1_3681(
      {stage115[39]},
      {stage115[177]}
   );
   gpc1_1 gpc1_1_3682(
      {stage115[40]},
      {stage115[178]}
   );
   gpc1_1 gpc1_1_3683(
      {stage115[41]},
      {stage115[179]}
   );
   gpc1_1 gpc1_1_3684(
      {stage115[42]},
      {stage115[180]}
   );
   gpc1_1 gpc1_1_3685(
      {stage115[43]},
      {stage115[181]}
   );
   gpc606_5 gpc606_5_3686(
      {stage115[44], stage115[45], stage115[46], stage115[47], stage115[48], stage115[49]},
      {stage117[0], stage117[1], stage117[2], stage117[3], stage117[4], stage117[5]},
      {stage119[128], stage118[132], stage117[145], stage116[152], stage115[182]}
   );
   gpc606_5 gpc606_5_3687(
      {stage115[50], stage115[51], stage115[52], stage115[53], stage115[54], stage115[55]},
      {stage117[6], stage117[7], stage117[8], stage117[9], stage117[10], stage117[11]},
      {stage119[129], stage118[133], stage117[146], stage116[153], stage115[183]}
   );
   gpc606_5 gpc606_5_3688(
      {stage115[56], stage115[57], stage115[58], stage115[59], stage115[60], stage115[61]},
      {stage117[12], stage117[13], stage117[14], stage117[15], stage117[16], stage117[17]},
      {stage119[130], stage118[134], stage117[147], stage116[154], stage115[184]}
   );
   gpc606_5 gpc606_5_3689(
      {stage115[62], stage115[63], stage115[64], stage115[65], stage115[66], stage115[67]},
      {stage117[18], stage117[19], stage117[20], stage117[21], stage117[22], stage117[23]},
      {stage119[131], stage118[135], stage117[148], stage116[155], stage115[185]}
   );
   gpc606_5 gpc606_5_3690(
      {stage115[68], stage115[69], stage115[70], stage115[71], stage115[72], stage115[73]},
      {stage117[24], stage117[25], stage117[26], stage117[27], stage117[28], stage117[29]},
      {stage119[132], stage118[136], stage117[149], stage116[156], stage115[186]}
   );
   gpc606_5 gpc606_5_3691(
      {stage115[74], stage115[75], stage115[76], stage115[77], stage115[78], stage115[79]},
      {stage117[30], stage117[31], stage117[32], stage117[33], stage117[34], stage117[35]},
      {stage119[133], stage118[137], stage117[150], stage116[157], stage115[187]}
   );
   gpc606_5 gpc606_5_3692(
      {stage115[80], stage115[81], stage115[82], stage115[83], stage115[84], stage115[85]},
      {stage117[36], stage117[37], stage117[38], stage117[39], stage117[40], stage117[41]},
      {stage119[134], stage118[138], stage117[151], stage116[158], stage115[188]}
   );
   gpc606_5 gpc606_5_3693(
      {stage115[86], stage115[87], stage115[88], stage115[89], stage115[90], stage115[91]},
      {stage117[42], stage117[43], stage117[44], stage117[45], stage117[46], stage117[47]},
      {stage119[135], stage118[139], stage117[152], stage116[159], stage115[189]}
   );
   gpc606_5 gpc606_5_3694(
      {stage115[92], stage115[93], stage115[94], stage115[95], stage115[96], stage115[97]},
      {stage117[48], stage117[49], stage117[50], stage117[51], stage117[52], stage117[53]},
      {stage119[136], stage118[140], stage117[153], stage116[160], stage115[190]}
   );
   gpc606_5 gpc606_5_3695(
      {stage115[98], stage115[99], stage115[100], stage115[101], stage115[102], stage115[103]},
      {stage117[54], stage117[55], stage117[56], stage117[57], stage117[58], stage117[59]},
      {stage119[137], stage118[141], stage117[154], stage116[161], stage115[191]}
   );
   gpc606_5 gpc606_5_3696(
      {stage115[104], stage115[105], stage115[106], stage115[107], stage115[108], stage115[109]},
      {stage117[60], stage117[61], stage117[62], stage117[63], stage117[64], stage117[65]},
      {stage119[138], stage118[142], stage117[155], stage116[162], stage115[192]}
   );
   gpc606_5 gpc606_5_3697(
      {stage115[110], stage115[111], stage115[112], stage115[113], stage115[114], stage115[115]},
      {stage117[66], stage117[67], stage117[68], stage117[69], stage117[70], stage117[71]},
      {stage119[139], stage118[143], stage117[156], stage116[163], stage115[193]}
   );
   gpc606_5 gpc606_5_3698(
      {stage115[116], stage115[117], stage115[118], stage115[119], stage115[120], stage115[121]},
      {stage117[72], stage117[73], stage117[74], stage117[75], stage117[76], stage117[77]},
      {stage119[140], stage118[144], stage117[157], stage116[164], stage115[194]}
   );
   gpc606_5 gpc606_5_3699(
      {stage115[122], stage115[123], stage115[124], stage115[125], stage115[126], stage115[127]},
      {stage117[78], stage117[79], stage117[80], stage117[81], stage117[82], stage117[83]},
      {stage119[141], stage118[145], stage117[158], stage116[165], stage115[195]}
   );
   gpc1_1 gpc1_1_3700(
      {stage116[42]},
      {stage116[166]}
   );
   gpc1_1 gpc1_1_3701(
      {stage116[43]},
      {stage116[167]}
   );
   gpc1_1 gpc1_1_3702(
      {stage116[44]},
      {stage116[168]}
   );
   gpc1_1 gpc1_1_3703(
      {stage116[45]},
      {stage116[169]}
   );
   gpc1_1 gpc1_1_3704(
      {stage116[46]},
      {stage116[170]}
   );
   gpc1_1 gpc1_1_3705(
      {stage116[47]},
      {stage116[171]}
   );
   gpc1_1 gpc1_1_3706(
      {stage116[48]},
      {stage116[172]}
   );
   gpc1_1 gpc1_1_3707(
      {stage116[49]},
      {stage116[173]}
   );
   gpc606_5 gpc606_5_3708(
      {stage116[50], stage116[51], stage116[52], stage116[53], stage116[54], stage116[55]},
      {stage118[0], stage118[1], stage118[2], stage118[3], stage118[4], stage118[5]},
      {stage120[128], stage119[142], stage118[146], stage117[159], stage116[174]}
   );
   gpc606_5 gpc606_5_3709(
      {stage116[56], stage116[57], stage116[58], stage116[59], stage116[60], stage116[61]},
      {stage118[6], stage118[7], stage118[8], stage118[9], stage118[10], stage118[11]},
      {stage120[129], stage119[143], stage118[147], stage117[160], stage116[175]}
   );
   gpc606_5 gpc606_5_3710(
      {stage116[62], stage116[63], stage116[64], stage116[65], stage116[66], stage116[67]},
      {stage118[12], stage118[13], stage118[14], stage118[15], stage118[16], stage118[17]},
      {stage120[130], stage119[144], stage118[148], stage117[161], stage116[176]}
   );
   gpc606_5 gpc606_5_3711(
      {stage116[68], stage116[69], stage116[70], stage116[71], stage116[72], stage116[73]},
      {stage118[18], stage118[19], stage118[20], stage118[21], stage118[22], stage118[23]},
      {stage120[131], stage119[145], stage118[149], stage117[162], stage116[177]}
   );
   gpc606_5 gpc606_5_3712(
      {stage116[74], stage116[75], stage116[76], stage116[77], stage116[78], stage116[79]},
      {stage118[24], stage118[25], stage118[26], stage118[27], stage118[28], stage118[29]},
      {stage120[132], stage119[146], stage118[150], stage117[163], stage116[178]}
   );
   gpc606_5 gpc606_5_3713(
      {stage116[80], stage116[81], stage116[82], stage116[83], stage116[84], stage116[85]},
      {stage118[30], stage118[31], stage118[32], stage118[33], stage118[34], stage118[35]},
      {stage120[133], stage119[147], stage118[151], stage117[164], stage116[179]}
   );
   gpc606_5 gpc606_5_3714(
      {stage116[86], stage116[87], stage116[88], stage116[89], stage116[90], stage116[91]},
      {stage118[36], stage118[37], stage118[38], stage118[39], stage118[40], stage118[41]},
      {stage120[134], stage119[148], stage118[152], stage117[165], stage116[180]}
   );
   gpc606_5 gpc606_5_3715(
      {stage116[92], stage116[93], stage116[94], stage116[95], stage116[96], stage116[97]},
      {stage118[42], stage118[43], stage118[44], stage118[45], stage118[46], stage118[47]},
      {stage120[135], stage119[149], stage118[153], stage117[166], stage116[181]}
   );
   gpc606_5 gpc606_5_3716(
      {stage116[98], stage116[99], stage116[100], stage116[101], stage116[102], stage116[103]},
      {stage118[48], stage118[49], stage118[50], stage118[51], stage118[52], stage118[53]},
      {stage120[136], stage119[150], stage118[154], stage117[167], stage116[182]}
   );
   gpc606_5 gpc606_5_3717(
      {stage116[104], stage116[105], stage116[106], stage116[107], stage116[108], stage116[109]},
      {stage118[54], stage118[55], stage118[56], stage118[57], stage118[58], stage118[59]},
      {stage120[137], stage119[151], stage118[155], stage117[168], stage116[183]}
   );
   gpc606_5 gpc606_5_3718(
      {stage116[110], stage116[111], stage116[112], stage116[113], stage116[114], stage116[115]},
      {stage118[60], stage118[61], stage118[62], stage118[63], stage118[64], stage118[65]},
      {stage120[138], stage119[152], stage118[156], stage117[169], stage116[184]}
   );
   gpc606_5 gpc606_5_3719(
      {stage116[116], stage116[117], stage116[118], stage116[119], stage116[120], stage116[121]},
      {stage118[66], stage118[67], stage118[68], stage118[69], stage118[70], stage118[71]},
      {stage120[139], stage119[153], stage118[157], stage117[170], stage116[185]}
   );
   gpc606_5 gpc606_5_3720(
      {stage116[122], stage116[123], stage116[124], stage116[125], stage116[126], stage116[127]},
      {stage118[72], stage118[73], stage118[74], stage118[75], stage118[76], stage118[77]},
      {stage120[140], stage119[154], stage118[158], stage117[171], stage116[186]}
   );
   gpc1_1 gpc1_1_3721(
      {stage117[84]},
      {stage117[172]}
   );
   gpc1_1 gpc1_1_3722(
      {stage117[85]},
      {stage117[173]}
   );
   gpc1_1 gpc1_1_3723(
      {stage117[86]},
      {stage117[174]}
   );
   gpc1_1 gpc1_1_3724(
      {stage117[87]},
      {stage117[175]}
   );
   gpc1_1 gpc1_1_3725(
      {stage117[88]},
      {stage117[176]}
   );
   gpc1_1 gpc1_1_3726(
      {stage117[89]},
      {stage117[177]}
   );
   gpc1_1 gpc1_1_3727(
      {stage117[90]},
      {stage117[178]}
   );
   gpc1_1 gpc1_1_3728(
      {stage117[91]},
      {stage117[179]}
   );
   gpc1_1 gpc1_1_3729(
      {stage117[92]},
      {stage117[180]}
   );
   gpc1_1 gpc1_1_3730(
      {stage117[93]},
      {stage117[181]}
   );
   gpc1_1 gpc1_1_3731(
      {stage117[94]},
      {stage117[182]}
   );
   gpc1_1 gpc1_1_3732(
      {stage117[95]},
      {stage117[183]}
   );
   gpc1_1 gpc1_1_3733(
      {stage117[96]},
      {stage117[184]}
   );
   gpc1_1 gpc1_1_3734(
      {stage117[97]},
      {stage117[185]}
   );
   gpc1_1 gpc1_1_3735(
      {stage117[98]},
      {stage117[186]}
   );
   gpc1_1 gpc1_1_3736(
      {stage117[99]},
      {stage117[187]}
   );
   gpc1_1 gpc1_1_3737(
      {stage117[100]},
      {stage117[188]}
   );
   gpc1_1 gpc1_1_3738(
      {stage117[101]},
      {stage117[189]}
   );
   gpc1_1 gpc1_1_3739(
      {stage117[102]},
      {stage117[190]}
   );
   gpc1_1 gpc1_1_3740(
      {stage117[103]},
      {stage117[191]}
   );
   gpc606_5 gpc606_5_3741(
      {stage117[104], stage117[105], stage117[106], stage117[107], stage117[108], stage117[109]},
      {stage119[0], stage119[1], stage119[2], stage119[3], stage119[4], stage119[5]},
      {stage121[128], stage120[141], stage119[155], stage118[159], stage117[192]}
   );
   gpc606_5 gpc606_5_3742(
      {stage117[110], stage117[111], stage117[112], stage117[113], stage117[114], stage117[115]},
      {stage119[6], stage119[7], stage119[8], stage119[9], stage119[10], stage119[11]},
      {stage121[129], stage120[142], stage119[156], stage118[160], stage117[193]}
   );
   gpc606_5 gpc606_5_3743(
      {stage117[116], stage117[117], stage117[118], stage117[119], stage117[120], stage117[121]},
      {stage119[12], stage119[13], stage119[14], stage119[15], stage119[16], stage119[17]},
      {stage121[130], stage120[143], stage119[157], stage118[161], stage117[194]}
   );
   gpc606_5 gpc606_5_3744(
      {stage117[122], stage117[123], stage117[124], stage117[125], stage117[126], stage117[127]},
      {stage119[18], stage119[19], stage119[20], stage119[21], stage119[22], stage119[23]},
      {stage121[131], stage120[144], stage119[158], stage118[162], stage117[195]}
   );
   gpc1_1 gpc1_1_3745(
      {stage118[78]},
      {stage118[163]}
   );
   gpc1_1 gpc1_1_3746(
      {stage118[79]},
      {stage118[164]}
   );
   gpc1_1 gpc1_1_3747(
      {stage118[80]},
      {stage118[165]}
   );
   gpc1_1 gpc1_1_3748(
      {stage118[81]},
      {stage118[166]}
   );
   gpc1_1 gpc1_1_3749(
      {stage118[82]},
      {stage118[167]}
   );
   gpc1_1 gpc1_1_3750(
      {stage118[83]},
      {stage118[168]}
   );
   gpc1_1 gpc1_1_3751(
      {stage118[84]},
      {stage118[169]}
   );
   gpc1_1 gpc1_1_3752(
      {stage118[85]},
      {stage118[170]}
   );
   gpc1_1 gpc1_1_3753(
      {stage118[86]},
      {stage118[171]}
   );
   gpc1_1 gpc1_1_3754(
      {stage118[87]},
      {stage118[172]}
   );
   gpc1_1 gpc1_1_3755(
      {stage118[88]},
      {stage118[173]}
   );
   gpc1_1 gpc1_1_3756(
      {stage118[89]},
      {stage118[174]}
   );
   gpc1_1 gpc1_1_3757(
      {stage118[90]},
      {stage118[175]}
   );
   gpc1_1 gpc1_1_3758(
      {stage118[91]},
      {stage118[176]}
   );
   gpc606_5 gpc606_5_3759(
      {stage118[92], stage118[93], stage118[94], stage118[95], stage118[96], stage118[97]},
      {stage120[0], stage120[1], stage120[2], stage120[3], stage120[4], stage120[5]},
      {stage122[128], stage121[132], stage120[145], stage119[159], stage118[177]}
   );
   gpc606_5 gpc606_5_3760(
      {stage118[98], stage118[99], stage118[100], stage118[101], stage118[102], stage118[103]},
      {stage120[6], stage120[7], stage120[8], stage120[9], stage120[10], stage120[11]},
      {stage122[129], stage121[133], stage120[146], stage119[160], stage118[178]}
   );
   gpc606_5 gpc606_5_3761(
      {stage118[104], stage118[105], stage118[106], stage118[107], stage118[108], stage118[109]},
      {stage120[12], stage120[13], stage120[14], stage120[15], stage120[16], stage120[17]},
      {stage122[130], stage121[134], stage120[147], stage119[161], stage118[179]}
   );
   gpc606_5 gpc606_5_3762(
      {stage118[110], stage118[111], stage118[112], stage118[113], stage118[114], stage118[115]},
      {stage120[18], stage120[19], stage120[20], stage120[21], stage120[22], stage120[23]},
      {stage122[131], stage121[135], stage120[148], stage119[162], stage118[180]}
   );
   gpc606_5 gpc606_5_3763(
      {stage118[116], stage118[117], stage118[118], stage118[119], stage118[120], stage118[121]},
      {stage120[24], stage120[25], stage120[26], stage120[27], stage120[28], stage120[29]},
      {stage122[132], stage121[136], stage120[149], stage119[163], stage118[181]}
   );
   gpc606_5 gpc606_5_3764(
      {stage118[122], stage118[123], stage118[124], stage118[125], stage118[126], stage118[127]},
      {stage120[30], stage120[31], stage120[32], stage120[33], stage120[34], stage120[35]},
      {stage122[133], stage121[137], stage120[150], stage119[164], stage118[182]}
   );
   gpc1_1 gpc1_1_3765(
      {stage119[24]},
      {stage119[165]}
   );
   gpc1_1 gpc1_1_3766(
      {stage119[25]},
      {stage119[166]}
   );
   gpc606_5 gpc606_5_3767(
      {stage119[26], stage119[27], stage119[28], stage119[29], stage119[30], stage119[31]},
      {stage121[0], stage121[1], stage121[2], stage121[3], stage121[4], stage121[5]},
      {stage123[128], stage122[134], stage121[138], stage120[151], stage119[167]}
   );
   gpc606_5 gpc606_5_3768(
      {stage119[32], stage119[33], stage119[34], stage119[35], stage119[36], stage119[37]},
      {stage121[6], stage121[7], stage121[8], stage121[9], stage121[10], stage121[11]},
      {stage123[129], stage122[135], stage121[139], stage120[152], stage119[168]}
   );
   gpc606_5 gpc606_5_3769(
      {stage119[38], stage119[39], stage119[40], stage119[41], stage119[42], stage119[43]},
      {stage121[12], stage121[13], stage121[14], stage121[15], stage121[16], stage121[17]},
      {stage123[130], stage122[136], stage121[140], stage120[153], stage119[169]}
   );
   gpc606_5 gpc606_5_3770(
      {stage119[44], stage119[45], stage119[46], stage119[47], stage119[48], stage119[49]},
      {stage121[18], stage121[19], stage121[20], stage121[21], stage121[22], stage121[23]},
      {stage123[131], stage122[137], stage121[141], stage120[154], stage119[170]}
   );
   gpc606_5 gpc606_5_3771(
      {stage119[50], stage119[51], stage119[52], stage119[53], stage119[54], stage119[55]},
      {stage121[24], stage121[25], stage121[26], stage121[27], stage121[28], stage121[29]},
      {stage123[132], stage122[138], stage121[142], stage120[155], stage119[171]}
   );
   gpc606_5 gpc606_5_3772(
      {stage119[56], stage119[57], stage119[58], stage119[59], stage119[60], stage119[61]},
      {stage121[30], stage121[31], stage121[32], stage121[33], stage121[34], stage121[35]},
      {stage123[133], stage122[139], stage121[143], stage120[156], stage119[172]}
   );
   gpc606_5 gpc606_5_3773(
      {stage119[62], stage119[63], stage119[64], stage119[65], stage119[66], stage119[67]},
      {stage121[36], stage121[37], stage121[38], stage121[39], stage121[40], stage121[41]},
      {stage123[134], stage122[140], stage121[144], stage120[157], stage119[173]}
   );
   gpc606_5 gpc606_5_3774(
      {stage119[68], stage119[69], stage119[70], stage119[71], stage119[72], stage119[73]},
      {stage121[42], stage121[43], stage121[44], stage121[45], stage121[46], stage121[47]},
      {stage123[135], stage122[141], stage121[145], stage120[158], stage119[174]}
   );
   gpc606_5 gpc606_5_3775(
      {stage119[74], stage119[75], stage119[76], stage119[77], stage119[78], stage119[79]},
      {stage121[48], stage121[49], stage121[50], stage121[51], stage121[52], stage121[53]},
      {stage123[136], stage122[142], stage121[146], stage120[159], stage119[175]}
   );
   gpc606_5 gpc606_5_3776(
      {stage119[80], stage119[81], stage119[82], stage119[83], stage119[84], stage119[85]},
      {stage121[54], stage121[55], stage121[56], stage121[57], stage121[58], stage121[59]},
      {stage123[137], stage122[143], stage121[147], stage120[160], stage119[176]}
   );
   gpc606_5 gpc606_5_3777(
      {stage119[86], stage119[87], stage119[88], stage119[89], stage119[90], stage119[91]},
      {stage121[60], stage121[61], stage121[62], stage121[63], stage121[64], stage121[65]},
      {stage123[138], stage122[144], stage121[148], stage120[161], stage119[177]}
   );
   gpc606_5 gpc606_5_3778(
      {stage119[92], stage119[93], stage119[94], stage119[95], stage119[96], stage119[97]},
      {stage121[66], stage121[67], stage121[68], stage121[69], stage121[70], stage121[71]},
      {stage123[139], stage122[145], stage121[149], stage120[162], stage119[178]}
   );
   gpc606_5 gpc606_5_3779(
      {stage119[98], stage119[99], stage119[100], stage119[101], stage119[102], stage119[103]},
      {stage121[72], stage121[73], stage121[74], stage121[75], stage121[76], stage121[77]},
      {stage123[140], stage122[146], stage121[150], stage120[163], stage119[179]}
   );
   gpc606_5 gpc606_5_3780(
      {stage119[104], stage119[105], stage119[106], stage119[107], stage119[108], stage119[109]},
      {stage121[78], stage121[79], stage121[80], stage121[81], stage121[82], stage121[83]},
      {stage123[141], stage122[147], stage121[151], stage120[164], stage119[180]}
   );
   gpc606_5 gpc606_5_3781(
      {stage119[110], stage119[111], stage119[112], stage119[113], stage119[114], stage119[115]},
      {stage121[84], stage121[85], stage121[86], stage121[87], stage121[88], stage121[89]},
      {stage123[142], stage122[148], stage121[152], stage120[165], stage119[181]}
   );
   gpc606_5 gpc606_5_3782(
      {stage119[116], stage119[117], stage119[118], stage119[119], stage119[120], stage119[121]},
      {stage121[90], stage121[91], stage121[92], stage121[93], stage121[94], stage121[95]},
      {stage123[143], stage122[149], stage121[153], stage120[166], stage119[182]}
   );
   gpc606_5 gpc606_5_3783(
      {stage119[122], stage119[123], stage119[124], stage119[125], stage119[126], stage119[127]},
      {stage121[96], stage121[97], stage121[98], stage121[99], stage121[100], stage121[101]},
      {stage123[144], stage122[150], stage121[154], stage120[167], stage119[183]}
   );
   gpc1_1 gpc1_1_3784(
      {stage120[36]},
      {stage120[168]}
   );
   gpc1_1 gpc1_1_3785(
      {stage120[37]},
      {stage120[169]}
   );
   gpc606_5 gpc606_5_3786(
      {stage120[38], stage120[39], stage120[40], stage120[41], stage120[42], stage120[43]},
      {stage122[0], stage122[1], stage122[2], stage122[3], stage122[4], stage122[5]},
      {stage124[128], stage123[145], stage122[151], stage121[155], stage120[170]}
   );
   gpc606_5 gpc606_5_3787(
      {stage120[44], stage120[45], stage120[46], stage120[47], stage120[48], stage120[49]},
      {stage122[6], stage122[7], stage122[8], stage122[9], stage122[10], stage122[11]},
      {stage124[129], stage123[146], stage122[152], stage121[156], stage120[171]}
   );
   gpc606_5 gpc606_5_3788(
      {stage120[50], stage120[51], stage120[52], stage120[53], stage120[54], stage120[55]},
      {stage122[12], stage122[13], stage122[14], stage122[15], stage122[16], stage122[17]},
      {stage124[130], stage123[147], stage122[153], stage121[157], stage120[172]}
   );
   gpc606_5 gpc606_5_3789(
      {stage120[56], stage120[57], stage120[58], stage120[59], stage120[60], stage120[61]},
      {stage122[18], stage122[19], stage122[20], stage122[21], stage122[22], stage122[23]},
      {stage124[131], stage123[148], stage122[154], stage121[158], stage120[173]}
   );
   gpc606_5 gpc606_5_3790(
      {stage120[62], stage120[63], stage120[64], stage120[65], stage120[66], stage120[67]},
      {stage122[24], stage122[25], stage122[26], stage122[27], stage122[28], stage122[29]},
      {stage124[132], stage123[149], stage122[155], stage121[159], stage120[174]}
   );
   gpc606_5 gpc606_5_3791(
      {stage120[68], stage120[69], stage120[70], stage120[71], stage120[72], stage120[73]},
      {stage122[30], stage122[31], stage122[32], stage122[33], stage122[34], stage122[35]},
      {stage124[133], stage123[150], stage122[156], stage121[160], stage120[175]}
   );
   gpc606_5 gpc606_5_3792(
      {stage120[74], stage120[75], stage120[76], stage120[77], stage120[78], stage120[79]},
      {stage122[36], stage122[37], stage122[38], stage122[39], stage122[40], stage122[41]},
      {stage124[134], stage123[151], stage122[157], stage121[161], stage120[176]}
   );
   gpc606_5 gpc606_5_3793(
      {stage120[80], stage120[81], stage120[82], stage120[83], stage120[84], stage120[85]},
      {stage122[42], stage122[43], stage122[44], stage122[45], stage122[46], stage122[47]},
      {stage124[135], stage123[152], stage122[158], stage121[162], stage120[177]}
   );
   gpc606_5 gpc606_5_3794(
      {stage120[86], stage120[87], stage120[88], stage120[89], stage120[90], stage120[91]},
      {stage122[48], stage122[49], stage122[50], stage122[51], stage122[52], stage122[53]},
      {stage124[136], stage123[153], stage122[159], stage121[163], stage120[178]}
   );
   gpc606_5 gpc606_5_3795(
      {stage120[92], stage120[93], stage120[94], stage120[95], stage120[96], stage120[97]},
      {stage122[54], stage122[55], stage122[56], stage122[57], stage122[58], stage122[59]},
      {stage124[137], stage123[154], stage122[160], stage121[164], stage120[179]}
   );
   gpc606_5 gpc606_5_3796(
      {stage120[98], stage120[99], stage120[100], stage120[101], stage120[102], stage120[103]},
      {stage122[60], stage122[61], stage122[62], stage122[63], stage122[64], stage122[65]},
      {stage124[138], stage123[155], stage122[161], stage121[165], stage120[180]}
   );
   gpc606_5 gpc606_5_3797(
      {stage120[104], stage120[105], stage120[106], stage120[107], stage120[108], stage120[109]},
      {stage122[66], stage122[67], stage122[68], stage122[69], stage122[70], stage122[71]},
      {stage124[139], stage123[156], stage122[162], stage121[166], stage120[181]}
   );
   gpc606_5 gpc606_5_3798(
      {stage120[110], stage120[111], stage120[112], stage120[113], stage120[114], stage120[115]},
      {stage122[72], stage122[73], stage122[74], stage122[75], stage122[76], stage122[77]},
      {stage124[140], stage123[157], stage122[163], stage121[167], stage120[182]}
   );
   gpc606_5 gpc606_5_3799(
      {stage120[116], stage120[117], stage120[118], stage120[119], stage120[120], stage120[121]},
      {stage122[78], stage122[79], stage122[80], stage122[81], stage122[82], stage122[83]},
      {stage124[141], stage123[158], stage122[164], stage121[168], stage120[183]}
   );
   gpc606_5 gpc606_5_3800(
      {stage120[122], stage120[123], stage120[124], stage120[125], stage120[126], stage120[127]},
      {stage122[84], stage122[85], stage122[86], stage122[87], stage122[88], stage122[89]},
      {stage124[142], stage123[159], stage122[165], stage121[169], stage120[184]}
   );
   gpc1_1 gpc1_1_3801(
      {stage121[102]},
      {stage121[170]}
   );
   gpc1_1 gpc1_1_3802(
      {stage121[103]},
      {stage121[171]}
   );
   gpc606_5 gpc606_5_3803(
      {stage121[104], stage121[105], stage121[106], stage121[107], stage121[108], stage121[109]},
      {stage123[0], stage123[1], stage123[2], stage123[3], stage123[4], stage123[5]},
      {stage125[128], stage124[143], stage123[160], stage122[166], stage121[172]}
   );
   gpc606_5 gpc606_5_3804(
      {stage121[110], stage121[111], stage121[112], stage121[113], stage121[114], stage121[115]},
      {stage123[6], stage123[7], stage123[8], stage123[9], stage123[10], stage123[11]},
      {stage125[129], stage124[144], stage123[161], stage122[167], stage121[173]}
   );
   gpc606_5 gpc606_5_3805(
      {stage121[116], stage121[117], stage121[118], stage121[119], stage121[120], stage121[121]},
      {stage123[12], stage123[13], stage123[14], stage123[15], stage123[16], stage123[17]},
      {stage125[130], stage124[145], stage123[162], stage122[168], stage121[174]}
   );
   gpc606_5 gpc606_5_3806(
      {stage121[122], stage121[123], stage121[124], stage121[125], stage121[126], stage121[127]},
      {stage123[18], stage123[19], stage123[20], stage123[21], stage123[22], stage123[23]},
      {stage125[131], stage124[146], stage123[163], stage122[169], stage121[175]}
   );
   gpc1_1 gpc1_1_3807(
      {stage122[90]},
      {stage122[170]}
   );
   gpc1_1 gpc1_1_3808(
      {stage122[91]},
      {stage122[171]}
   );
   gpc1_1 gpc1_1_3809(
      {stage122[92]},
      {stage122[172]}
   );
   gpc1_1 gpc1_1_3810(
      {stage122[93]},
      {stage122[173]}
   );
   gpc1_1 gpc1_1_3811(
      {stage122[94]},
      {stage122[174]}
   );
   gpc1_1 gpc1_1_3812(
      {stage122[95]},
      {stage122[175]}
   );
   gpc1_1 gpc1_1_3813(
      {stage122[96]},
      {stage122[176]}
   );
   gpc1_1 gpc1_1_3814(
      {stage122[97]},
      {stage122[177]}
   );
   gpc1_1 gpc1_1_3815(
      {stage122[98]},
      {stage122[178]}
   );
   gpc1_1 gpc1_1_3816(
      {stage122[99]},
      {stage122[179]}
   );
   gpc1_1 gpc1_1_3817(
      {stage122[100]},
      {stage122[180]}
   );
   gpc1_1 gpc1_1_3818(
      {stage122[101]},
      {stage122[181]}
   );
   gpc606_5 gpc606_5_3819(
      {stage122[102], stage122[103], stage122[104], stage122[105], stage122[106], stage122[107]},
      {stage124[0], stage124[1], stage124[2], stage124[3], stage124[4], stage124[5]},
      {stage126[128], stage125[132], stage124[147], stage123[164], stage122[182]}
   );
   gpc2135_5 gpc2135_5_3820(
      {stage122[108], stage122[109], stage122[110], stage122[111], stage122[112]},
      {stage123[24], stage123[25], stage123[26]},
      {stage124[6]},
      {stage125[0], stage125[1]},
      {stage126[129], stage125[133], stage124[148], stage123[165], stage122[183]}
   );
   gpc2135_5 gpc2135_5_3821(
      {stage122[113], stage122[114], stage122[115], stage122[116], stage122[117]},
      {stage123[27], stage123[28], stage123[29]},
      {stage124[7]},
      {stage125[2], stage125[3]},
      {stage126[130], stage125[134], stage124[149], stage123[166], stage122[184]}
   );
   gpc2135_5 gpc2135_5_3822(
      {stage122[118], stage122[119], stage122[120], stage122[121], stage122[122]},
      {stage123[30], stage123[31], stage123[32]},
      {stage124[8]},
      {stage125[4], stage125[5]},
      {stage126[131], stage125[135], stage124[150], stage123[167], stage122[185]}
   );
   gpc2135_5 gpc2135_5_3823(
      {stage122[123], stage122[124], stage122[125], stage122[126], stage122[127]},
      {stage123[33], stage123[34], stage123[35]},
      {stage124[9]},
      {stage125[6], stage125[7]},
      {stage126[132], stage125[136], stage124[151], stage123[168], stage122[186]}
   );
   gpc1_1 gpc1_1_3824(
      {stage123[36]},
      {stage123[169]}
   );
   gpc1_1 gpc1_1_3825(
      {stage123[37]},
      {stage123[170]}
   );
   gpc1_1 gpc1_1_3826(
      {stage123[38]},
      {stage123[171]}
   );
   gpc1_1 gpc1_1_3827(
      {stage123[39]},
      {stage123[172]}
   );
   gpc1_1 gpc1_1_3828(
      {stage123[40]},
      {stage123[173]}
   );
   gpc1_1 gpc1_1_3829(
      {stage123[41]},
      {stage123[174]}
   );
   gpc1_1 gpc1_1_3830(
      {stage123[42]},
      {stage123[175]}
   );
   gpc1_1 gpc1_1_3831(
      {stage123[43]},
      {stage123[176]}
   );
   gpc1_1 gpc1_1_3832(
      {stage123[44]},
      {stage123[177]}
   );
   gpc1_1 gpc1_1_3833(
      {stage123[45]},
      {stage123[178]}
   );
   gpc1_1 gpc1_1_3834(
      {stage123[46]},
      {stage123[179]}
   );
   gpc1_1 gpc1_1_3835(
      {stage123[47]},
      {stage123[180]}
   );
   gpc1_1 gpc1_1_3836(
      {stage123[48]},
      {stage123[181]}
   );
   gpc1_1 gpc1_1_3837(
      {stage123[49]},
      {stage123[182]}
   );
   gpc1_1 gpc1_1_3838(
      {stage123[50]},
      {stage123[183]}
   );
   gpc1_1 gpc1_1_3839(
      {stage123[51]},
      {stage123[184]}
   );
   gpc1_1 gpc1_1_3840(
      {stage123[52]},
      {stage123[185]}
   );
   gpc1_1 gpc1_1_3841(
      {stage123[53]},
      {stage123[186]}
   );
   gpc1_1 gpc1_1_3842(
      {stage123[54]},
      {stage123[187]}
   );
   gpc1_1 gpc1_1_3843(
      {stage123[55]},
      {stage123[188]}
   );
   gpc1_1 gpc1_1_3844(
      {stage123[56]},
      {stage123[189]}
   );
   gpc1_1 gpc1_1_3845(
      {stage123[57]},
      {stage123[190]}
   );
   gpc1_1 gpc1_1_3846(
      {stage123[58]},
      {stage123[191]}
   );
   gpc1_1 gpc1_1_3847(
      {stage123[59]},
      {stage123[192]}
   );
   gpc1_1 gpc1_1_3848(
      {stage123[60]},
      {stage123[193]}
   );
   gpc1_1 gpc1_1_3849(
      {stage123[61]},
      {stage123[194]}
   );
   gpc1_1 gpc1_1_3850(
      {stage123[62]},
      {stage123[195]}
   );
   gpc1_1 gpc1_1_3851(
      {stage123[63]},
      {stage123[196]}
   );
   gpc1_1 gpc1_1_3852(
      {stage123[64]},
      {stage123[197]}
   );
   gpc1_1 gpc1_1_3853(
      {stage123[65]},
      {stage123[198]}
   );
   gpc1_1 gpc1_1_3854(
      {stage123[66]},
      {stage123[199]}
   );
   gpc1_1 gpc1_1_3855(
      {stage123[67]},
      {stage123[200]}
   );
   gpc1_1 gpc1_1_3856(
      {stage123[68]},
      {stage123[201]}
   );
   gpc1_1 gpc1_1_3857(
      {stage123[69]},
      {stage123[202]}
   );
   gpc1_1 gpc1_1_3858(
      {stage123[70]},
      {stage123[203]}
   );
   gpc1_1 gpc1_1_3859(
      {stage123[71]},
      {stage123[204]}
   );
   gpc1_1 gpc1_1_3860(
      {stage123[72]},
      {stage123[205]}
   );
   gpc1_1 gpc1_1_3861(
      {stage123[73]},
      {stage123[206]}
   );
   gpc1_1 gpc1_1_3862(
      {stage123[74]},
      {stage123[207]}
   );
   gpc1_1 gpc1_1_3863(
      {stage123[75]},
      {stage123[208]}
   );
   gpc1_1 gpc1_1_3864(
      {stage123[76]},
      {stage123[209]}
   );
   gpc1_1 gpc1_1_3865(
      {stage123[77]},
      {stage123[210]}
   );
   gpc1_1 gpc1_1_3866(
      {stage123[78]},
      {stage123[211]}
   );
   gpc1_1 gpc1_1_3867(
      {stage123[79]},
      {stage123[212]}
   );
   gpc1_1 gpc1_1_3868(
      {stage123[80]},
      {stage123[213]}
   );
   gpc1_1 gpc1_1_3869(
      {stage123[81]},
      {stage123[214]}
   );
   gpc1_1 gpc1_1_3870(
      {stage123[82]},
      {stage123[215]}
   );
   gpc1_1 gpc1_1_3871(
      {stage123[83]},
      {stage123[216]}
   );
   gpc1_1 gpc1_1_3872(
      {stage123[84]},
      {stage123[217]}
   );
   gpc1_1 gpc1_1_3873(
      {stage123[85]},
      {stage123[218]}
   );
   gpc1_1 gpc1_1_3874(
      {stage123[86]},
      {stage123[219]}
   );
   gpc1_1 gpc1_1_3875(
      {stage123[87]},
      {stage123[220]}
   );
   gpc1_1 gpc1_1_3876(
      {stage123[88]},
      {stage123[221]}
   );
   gpc1_1 gpc1_1_3877(
      {stage123[89]},
      {stage123[222]}
   );
   gpc1_1 gpc1_1_3878(
      {stage123[90]},
      {stage123[223]}
   );
   gpc1_1 gpc1_1_3879(
      {stage123[91]},
      {stage123[224]}
   );
   gpc1_1 gpc1_1_3880(
      {stage123[92]},
      {stage123[225]}
   );
   gpc1_1 gpc1_1_3881(
      {stage123[93]},
      {stage123[226]}
   );
   gpc1_1 gpc1_1_3882(
      {stage123[94]},
      {stage123[227]}
   );
   gpc1_1 gpc1_1_3883(
      {stage123[95]},
      {stage123[228]}
   );
   gpc1_1 gpc1_1_3884(
      {stage123[96]},
      {stage123[229]}
   );
   gpc1_1 gpc1_1_3885(
      {stage123[97]},
      {stage123[230]}
   );
   gpc1_1 gpc1_1_3886(
      {stage123[98]},
      {stage123[231]}
   );
   gpc1_1 gpc1_1_3887(
      {stage123[99]},
      {stage123[232]}
   );
   gpc1_1 gpc1_1_3888(
      {stage123[100]},
      {stage123[233]}
   );
   gpc1_1 gpc1_1_3889(
      {stage123[101]},
      {stage123[234]}
   );
   gpc1_1 gpc1_1_3890(
      {stage123[102]},
      {stage123[235]}
   );
   gpc1_1 gpc1_1_3891(
      {stage123[103]},
      {stage123[236]}
   );
   gpc1_1 gpc1_1_3892(
      {stage123[104]},
      {stage123[237]}
   );
   gpc1_1 gpc1_1_3893(
      {stage123[105]},
      {stage123[238]}
   );
   gpc1_1 gpc1_1_3894(
      {stage123[106]},
      {stage123[239]}
   );
   gpc1_1 gpc1_1_3895(
      {stage123[107]},
      {stage123[240]}
   );
   gpc1_1 gpc1_1_3896(
      {stage123[108]},
      {stage123[241]}
   );
   gpc1_1 gpc1_1_3897(
      {stage123[109]},
      {stage123[242]}
   );
   gpc1_1 gpc1_1_3898(
      {stage123[110]},
      {stage123[243]}
   );
   gpc1_1 gpc1_1_3899(
      {stage123[111]},
      {stage123[244]}
   );
   gpc1_1 gpc1_1_3900(
      {stage123[112]},
      {stage123[245]}
   );
   gpc1_1 gpc1_1_3901(
      {stage123[113]},
      {stage123[246]}
   );
   gpc1_1 gpc1_1_3902(
      {stage123[114]},
      {stage123[247]}
   );
   gpc1_1 gpc1_1_3903(
      {stage123[115]},
      {stage123[248]}
   );
   gpc1_1 gpc1_1_3904(
      {stage123[116]},
      {stage123[249]}
   );
   gpc1_1 gpc1_1_3905(
      {stage123[117]},
      {stage123[250]}
   );
   gpc1_1 gpc1_1_3906(
      {stage123[118]},
      {stage123[251]}
   );
   gpc1_1 gpc1_1_3907(
      {stage123[119]},
      {stage123[252]}
   );
   gpc1_1 gpc1_1_3908(
      {stage123[120]},
      {stage123[253]}
   );
   gpc1_1 gpc1_1_3909(
      {stage123[121]},
      {stage123[254]}
   );
   gpc606_5 gpc606_5_3910(
      {stage123[122], stage123[123], stage123[124], stage123[125], stage123[126], stage123[127]},
      {stage125[8], stage125[9], stage125[10], stage125[11], stage125[12], stage125[13]},
      {stage127[128], stage126[133], stage125[137], stage124[152], stage123[255]}
   );
   gpc1_1 gpc1_1_3911(
      {stage124[10]},
      {stage124[153]}
   );
   gpc1_1 gpc1_1_3912(
      {stage124[11]},
      {stage124[154]}
   );
   gpc1_1 gpc1_1_3913(
      {stage124[12]},
      {stage124[155]}
   );
   gpc1_1 gpc1_1_3914(
      {stage124[13]},
      {stage124[156]}
   );
   gpc1_1 gpc1_1_3915(
      {stage124[14]},
      {stage124[157]}
   );
   gpc1_1 gpc1_1_3916(
      {stage124[15]},
      {stage124[158]}
   );
   gpc606_5 gpc606_5_3917(
      {stage124[16], stage124[17], stage124[18], stage124[19], stage124[20], stage124[21]},
      {stage126[0], stage126[1], stage126[2], stage126[3], stage126[4], stage126[5]},
      {stage128[0], stage127[129], stage126[134], stage125[138], stage124[159]}
   );
   gpc606_5 gpc606_5_3918(
      {stage124[22], stage124[23], stage124[24], stage124[25], stage124[26], stage124[27]},
      {stage126[6], stage126[7], stage126[8], stage126[9], stage126[10], stage126[11]},
      {stage128[1], stage127[130], stage126[135], stage125[139], stage124[160]}
   );
   gpc606_5 gpc606_5_3919(
      {stage124[28], stage124[29], stage124[30], stage124[31], stage124[32], stage124[33]},
      {stage126[12], stage126[13], stage126[14], stage126[15], stage126[16], stage126[17]},
      {stage128[2], stage127[131], stage126[136], stage125[140], stage124[161]}
   );
   gpc606_5 gpc606_5_3920(
      {stage124[34], stage124[35], stage124[36], stage124[37], stage124[38], stage124[39]},
      {stage126[18], stage126[19], stage126[20], stage126[21], stage126[22], stage126[23]},
      {stage128[3], stage127[132], stage126[137], stage125[141], stage124[162]}
   );
   gpc606_5 gpc606_5_3921(
      {stage124[40], stage124[41], stage124[42], stage124[43], stage124[44], stage124[45]},
      {stage126[24], stage126[25], stage126[26], stage126[27], stage126[28], stage126[29]},
      {stage128[4], stage127[133], stage126[138], stage125[142], stage124[163]}
   );
   gpc606_5 gpc606_5_3922(
      {stage124[46], stage124[47], stage124[48], stage124[49], stage124[50], stage124[51]},
      {stage126[30], stage126[31], stage126[32], stage126[33], stage126[34], stage126[35]},
      {stage128[5], stage127[134], stage126[139], stage125[143], stage124[164]}
   );
   gpc606_5 gpc606_5_3923(
      {stage124[52], stage124[53], stage124[54], stage124[55], stage124[56], stage124[57]},
      {stage126[36], stage126[37], stage126[38], stage126[39], stage126[40], stage126[41]},
      {stage128[6], stage127[135], stage126[140], stage125[144], stage124[165]}
   );
   gpc606_5 gpc606_5_3924(
      {stage124[58], stage124[59], stage124[60], stage124[61], stage124[62], stage124[63]},
      {stage126[42], stage126[43], stage126[44], stage126[45], stage126[46], stage126[47]},
      {stage128[7], stage127[136], stage126[141], stage125[145], stage124[166]}
   );
   gpc606_5 gpc606_5_3925(
      {stage124[64], stage124[65], stage124[66], stage124[67], stage124[68], stage124[69]},
      {stage126[48], stage126[49], stage126[50], stage126[51], stage126[52], stage126[53]},
      {stage128[8], stage127[137], stage126[142], stage125[146], stage124[167]}
   );
   gpc606_5 gpc606_5_3926(
      {stage124[70], stage124[71], stage124[72], stage124[73], stage124[74], stage124[75]},
      {stage126[54], stage126[55], stage126[56], stage126[57], stage126[58], stage126[59]},
      {stage128[9], stage127[138], stage126[143], stage125[147], stage124[168]}
   );
   gpc606_5 gpc606_5_3927(
      {stage124[76], stage124[77], stage124[78], stage124[79], stage124[80], stage124[81]},
      {stage126[60], stage126[61], stage126[62], stage126[63], stage126[64], stage126[65]},
      {stage128[10], stage127[139], stage126[144], stage125[148], stage124[169]}
   );
   gpc606_5 gpc606_5_3928(
      {stage124[82], stage124[83], stage124[84], stage124[85], stage124[86], stage124[87]},
      {stage126[66], stage126[67], stage126[68], stage126[69], stage126[70], stage126[71]},
      {stage128[11], stage127[140], stage126[145], stage125[149], stage124[170]}
   );
   gpc606_5 gpc606_5_3929(
      {stage124[88], stage124[89], stage124[90], stage124[91], stage124[92], stage124[93]},
      {stage126[72], stage126[73], stage126[74], stage126[75], stage126[76], stage126[77]},
      {stage128[12], stage127[141], stage126[146], stage125[150], stage124[171]}
   );
   gpc606_5 gpc606_5_3930(
      {stage124[94], stage124[95], stage124[96], stage124[97], stage124[98], stage124[99]},
      {stage126[78], stage126[79], stage126[80], stage126[81], stage126[82], stage126[83]},
      {stage128[13], stage127[142], stage126[147], stage125[151], stage124[172]}
   );
   gpc606_5 gpc606_5_3931(
      {stage124[100], stage124[101], stage124[102], stage124[103], stage124[104], stage124[105]},
      {stage126[84], stage126[85], stage126[86], stage126[87], stage126[88], stage126[89]},
      {stage128[14], stage127[143], stage126[148], stage125[152], stage124[173]}
   );
   gpc606_5 gpc606_5_3932(
      {stage124[106], stage124[107], stage124[108], stage124[109], stage124[110], stage124[111]},
      {stage126[90], stage126[91], stage126[92], stage126[93], stage126[94], stage126[95]},
      {stage128[15], stage127[144], stage126[149], stage125[153], stage124[174]}
   );
   gpc606_5 gpc606_5_3933(
      {stage124[112], stage124[113], stage124[114], stage124[115], stage124[116], stage124[117]},
      {stage126[96], stage126[97], stage126[98], stage126[99], stage126[100], stage126[101]},
      {stage128[16], stage127[145], stage126[150], stage125[154], stage124[175]}
   );
   gpc2135_5 gpc2135_5_3934(
      {stage124[118], stage124[119], stage124[120], stage124[121], stage124[122]},
      {stage125[14], stage125[15], stage125[16]},
      {stage126[102]},
      {stage127[0], stage127[1]},
      {stage128[17], stage127[146], stage126[151], stage125[155], stage124[176]}
   );
   gpc2135_5 gpc2135_5_3935(
      {stage124[123], stage124[124], stage124[125], stage124[126], stage124[127]},
      {stage125[17], stage125[18], stage125[19]},
      {stage126[103]},
      {stage127[2], stage127[3]},
      {stage128[18], stage127[147], stage126[152], stage125[156], stage124[177]}
   );
   gpc1_1 gpc1_1_3936(
      {stage125[20]},
      {stage125[157]}
   );
   gpc1_1 gpc1_1_3937(
      {stage125[21]},
      {stage125[158]}
   );
   gpc1_1 gpc1_1_3938(
      {stage125[22]},
      {stage125[159]}
   );
   gpc1_1 gpc1_1_3939(
      {stage125[23]},
      {stage125[160]}
   );
   gpc1_1 gpc1_1_3940(
      {stage125[24]},
      {stage125[161]}
   );
   gpc1_1 gpc1_1_3941(
      {stage125[25]},
      {stage125[162]}
   );
   gpc1_1 gpc1_1_3942(
      {stage125[26]},
      {stage125[163]}
   );
   gpc1_1 gpc1_1_3943(
      {stage125[27]},
      {stage125[164]}
   );
   gpc1_1 gpc1_1_3944(
      {stage125[28]},
      {stage125[165]}
   );
   gpc1_1 gpc1_1_3945(
      {stage125[29]},
      {stage125[166]}
   );
   gpc1_1 gpc1_1_3946(
      {stage125[30]},
      {stage125[167]}
   );
   gpc1_1 gpc1_1_3947(
      {stage125[31]},
      {stage125[168]}
   );
   gpc1_1 gpc1_1_3948(
      {stage125[32]},
      {stage125[169]}
   );
   gpc1_1 gpc1_1_3949(
      {stage125[33]},
      {stage125[170]}
   );
   gpc1_1 gpc1_1_3950(
      {stage125[34]},
      {stage125[171]}
   );
   gpc1_1 gpc1_1_3951(
      {stage125[35]},
      {stage125[172]}
   );
   gpc1_1 gpc1_1_3952(
      {stage125[36]},
      {stage125[173]}
   );
   gpc1_1 gpc1_1_3953(
      {stage125[37]},
      {stage125[174]}
   );
   gpc1_1 gpc1_1_3954(
      {stage125[38]},
      {stage125[175]}
   );
   gpc1_1 gpc1_1_3955(
      {stage125[39]},
      {stage125[176]}
   );
   gpc1_1 gpc1_1_3956(
      {stage125[40]},
      {stage125[177]}
   );
   gpc1_1 gpc1_1_3957(
      {stage125[41]},
      {stage125[178]}
   );
   gpc1_1 gpc1_1_3958(
      {stage125[42]},
      {stage125[179]}
   );
   gpc1_1 gpc1_1_3959(
      {stage125[43]},
      {stage125[180]}
   );
   gpc1_1 gpc1_1_3960(
      {stage125[44]},
      {stage125[181]}
   );
   gpc1_1 gpc1_1_3961(
      {stage125[45]},
      {stage125[182]}
   );
   gpc1_1 gpc1_1_3962(
      {stage125[46]},
      {stage125[183]}
   );
   gpc1_1 gpc1_1_3963(
      {stage125[47]},
      {stage125[184]}
   );
   gpc1_1 gpc1_1_3964(
      {stage125[48]},
      {stage125[185]}
   );
   gpc1_1 gpc1_1_3965(
      {stage125[49]},
      {stage125[186]}
   );
   gpc1_1 gpc1_1_3966(
      {stage125[50]},
      {stage125[187]}
   );
   gpc1_1 gpc1_1_3967(
      {stage125[51]},
      {stage125[188]}
   );
   gpc1_1 gpc1_1_3968(
      {stage125[52]},
      {stage125[189]}
   );
   gpc1_1 gpc1_1_3969(
      {stage125[53]},
      {stage125[190]}
   );
   gpc1_1 gpc1_1_3970(
      {stage125[54]},
      {stage125[191]}
   );
   gpc1_1 gpc1_1_3971(
      {stage125[55]},
      {stage125[192]}
   );
   gpc606_5 gpc606_5_3972(
      {stage125[56], stage125[57], stage125[58], stage125[59], stage125[60], stage125[61]},
      {stage127[4], stage127[5], stage127[6], stage127[7], stage127[8], stage127[9]},
      {stage129[0], stage128[19], stage127[148], stage126[153], stage125[193]}
   );
   gpc606_5 gpc606_5_3973(
      {stage125[62], stage125[63], stage125[64], stage125[65], stage125[66], stage125[67]},
      {stage127[10], stage127[11], stage127[12], stage127[13], stage127[14], stage127[15]},
      {stage129[1], stage128[20], stage127[149], stage126[154], stage125[194]}
   );
   gpc606_5 gpc606_5_3974(
      {stage125[68], stage125[69], stage125[70], stage125[71], stage125[72], stage125[73]},
      {stage127[16], stage127[17], stage127[18], stage127[19], stage127[20], stage127[21]},
      {stage129[2], stage128[21], stage127[150], stage126[155], stage125[195]}
   );
   gpc606_5 gpc606_5_3975(
      {stage125[74], stage125[75], stage125[76], stage125[77], stage125[78], stage125[79]},
      {stage127[22], stage127[23], stage127[24], stage127[25], stage127[26], stage127[27]},
      {stage129[3], stage128[22], stage127[151], stage126[156], stage125[196]}
   );
   gpc606_5 gpc606_5_3976(
      {stage125[80], stage125[81], stage125[82], stage125[83], stage125[84], stage125[85]},
      {stage127[28], stage127[29], stage127[30], stage127[31], stage127[32], stage127[33]},
      {stage129[4], stage128[23], stage127[152], stage126[157], stage125[197]}
   );
   gpc606_5 gpc606_5_3977(
      {stage125[86], stage125[87], stage125[88], stage125[89], stage125[90], stage125[91]},
      {stage127[34], stage127[35], stage127[36], stage127[37], stage127[38], stage127[39]},
      {stage129[5], stage128[24], stage127[153], stage126[158], stage125[198]}
   );
   gpc606_5 gpc606_5_3978(
      {stage125[92], stage125[93], stage125[94], stage125[95], stage125[96], stage125[97]},
      {stage127[40], stage127[41], stage127[42], stage127[43], stage127[44], stage127[45]},
      {stage129[6], stage128[25], stage127[154], stage126[159], stage125[199]}
   );
   gpc606_5 gpc606_5_3979(
      {stage125[98], stage125[99], stage125[100], stage125[101], stage125[102], stage125[103]},
      {stage127[46], stage127[47], stage127[48], stage127[49], stage127[50], stage127[51]},
      {stage129[7], stage128[26], stage127[155], stage126[160], stage125[200]}
   );
   gpc606_5 gpc606_5_3980(
      {stage125[104], stage125[105], stage125[106], stage125[107], stage125[108], stage125[109]},
      {stage127[52], stage127[53], stage127[54], stage127[55], stage127[56], stage127[57]},
      {stage129[8], stage128[27], stage127[156], stage126[161], stage125[201]}
   );
   gpc606_5 gpc606_5_3981(
      {stage125[110], stage125[111], stage125[112], stage125[113], stage125[114], stage125[115]},
      {stage127[58], stage127[59], stage127[60], stage127[61], stage127[62], stage127[63]},
      {stage129[9], stage128[28], stage127[157], stage126[162], stage125[202]}
   );
   gpc606_5 gpc606_5_3982(
      {stage125[116], stage125[117], stage125[118], stage125[119], stage125[120], stage125[121]},
      {stage127[64], stage127[65], stage127[66], stage127[67], stage127[68], stage127[69]},
      {stage129[10], stage128[29], stage127[158], stage126[163], stage125[203]}
   );
   gpc606_5 gpc606_5_3983(
      {stage125[122], stage125[123], stage125[124], stage125[125], stage125[126], stage125[127]},
      {stage127[70], stage127[71], stage127[72], stage127[73], stage127[74], stage127[75]},
      {stage129[11], stage128[30], stage127[159], stage126[164], stage125[204]}
   );
   gpc1_1 gpc1_1_3984(
      {stage126[104]},
      {stage126[165]}
   );
   gpc1_1 gpc1_1_3985(
      {stage126[105]},
      {stage126[166]}
   );
   gpc1_1 gpc1_1_3986(
      {stage126[106]},
      {stage126[167]}
   );
   gpc1_1 gpc1_1_3987(
      {stage126[107]},
      {stage126[168]}
   );
   gpc1_1 gpc1_1_3988(
      {stage126[108]},
      {stage126[169]}
   );
   gpc1_1 gpc1_1_3989(
      {stage126[109]},
      {stage126[170]}
   );
   gpc1_1 gpc1_1_3990(
      {stage126[110]},
      {stage126[171]}
   );
   gpc1_1 gpc1_1_3991(
      {stage126[111]},
      {stage126[172]}
   );
   gpc1_1 gpc1_1_3992(
      {stage126[112]},
      {stage126[173]}
   );
   gpc1_1 gpc1_1_3993(
      {stage126[113]},
      {stage126[174]}
   );
   gpc1_1 gpc1_1_3994(
      {stage126[114]},
      {stage126[175]}
   );
   gpc1_1 gpc1_1_3995(
      {stage126[115]},
      {stage126[176]}
   );
   gpc1_1 gpc1_1_3996(
      {stage126[116]},
      {stage126[177]}
   );
   gpc1_1 gpc1_1_3997(
      {stage126[117]},
      {stage126[178]}
   );
   gpc1_1 gpc1_1_3998(
      {stage126[118]},
      {stage126[179]}
   );
   gpc1_1 gpc1_1_3999(
      {stage126[119]},
      {stage126[180]}
   );
   gpc1_1 gpc1_1_4000(
      {stage126[120]},
      {stage126[181]}
   );
   gpc1_1 gpc1_1_4001(
      {stage126[121]},
      {stage126[182]}
   );
   gpc1_1 gpc1_1_4002(
      {stage126[122]},
      {stage126[183]}
   );
   gpc1_1 gpc1_1_4003(
      {stage126[123]},
      {stage126[184]}
   );
   gpc1_1 gpc1_1_4004(
      {stage126[124]},
      {stage126[185]}
   );
   gpc1_1 gpc1_1_4005(
      {stage126[125]},
      {stage126[186]}
   );
   gpc1_1 gpc1_1_4006(
      {stage126[126]},
      {stage126[187]}
   );
   gpc1_1 gpc1_1_4007(
      {stage126[127]},
      {stage126[188]}
   );
   gpc1_1 gpc1_1_4008(
      {stage127[76]},
      {stage127[160]}
   );
   gpc1_1 gpc1_1_4009(
      {stage127[77]},
      {stage127[161]}
   );
   gpc1_1 gpc1_1_4010(
      {stage127[78]},
      {stage127[162]}
   );
   gpc1_1 gpc1_1_4011(
      {stage127[79]},
      {stage127[163]}
   );
   gpc1_1 gpc1_1_4012(
      {stage127[80]},
      {stage127[164]}
   );
   gpc1_1 gpc1_1_4013(
      {stage127[81]},
      {stage127[165]}
   );
   gpc1_1 gpc1_1_4014(
      {stage127[82]},
      {stage127[166]}
   );
   gpc1_1 gpc1_1_4015(
      {stage127[83]},
      {stage127[167]}
   );
   gpc1_1 gpc1_1_4016(
      {stage127[84]},
      {stage127[168]}
   );
   gpc1_1 gpc1_1_4017(
      {stage127[85]},
      {stage127[169]}
   );
   gpc1_1 gpc1_1_4018(
      {stage127[86]},
      {stage127[170]}
   );
   gpc1_1 gpc1_1_4019(
      {stage127[87]},
      {stage127[171]}
   );
   gpc1_1 gpc1_1_4020(
      {stage127[88]},
      {stage127[172]}
   );
   gpc1_1 gpc1_1_4021(
      {stage127[89]},
      {stage127[173]}
   );
   gpc1_1 gpc1_1_4022(
      {stage127[90]},
      {stage127[174]}
   );
   gpc1_1 gpc1_1_4023(
      {stage127[91]},
      {stage127[175]}
   );
   gpc1_1 gpc1_1_4024(
      {stage127[92]},
      {stage127[176]}
   );
   gpc1_1 gpc1_1_4025(
      {stage127[93]},
      {stage127[177]}
   );
   gpc1_1 gpc1_1_4026(
      {stage127[94]},
      {stage127[178]}
   );
   gpc1_1 gpc1_1_4027(
      {stage127[95]},
      {stage127[179]}
   );
   gpc1_1 gpc1_1_4028(
      {stage127[96]},
      {stage127[180]}
   );
   gpc1_1 gpc1_1_4029(
      {stage127[97]},
      {stage127[181]}
   );
   gpc1_1 gpc1_1_4030(
      {stage127[98]},
      {stage127[182]}
   );
   gpc1_1 gpc1_1_4031(
      {stage127[99]},
      {stage127[183]}
   );
   gpc1_1 gpc1_1_4032(
      {stage127[100]},
      {stage127[184]}
   );
   gpc1_1 gpc1_1_4033(
      {stage127[101]},
      {stage127[185]}
   );
   gpc1_1 gpc1_1_4034(
      {stage127[102]},
      {stage127[186]}
   );
   gpc1_1 gpc1_1_4035(
      {stage127[103]},
      {stage127[187]}
   );
   gpc1_1 gpc1_1_4036(
      {stage127[104]},
      {stage127[188]}
   );
   gpc1_1 gpc1_1_4037(
      {stage127[105]},
      {stage127[189]}
   );
   gpc1_1 gpc1_1_4038(
      {stage127[106]},
      {stage127[190]}
   );
   gpc1_1 gpc1_1_4039(
      {stage127[107]},
      {stage127[191]}
   );
   gpc1_1 gpc1_1_4040(
      {stage127[108]},
      {stage127[192]}
   );
   gpc1_1 gpc1_1_4041(
      {stage127[109]},
      {stage127[193]}
   );
   gpc1_1 gpc1_1_4042(
      {stage127[110]},
      {stage127[194]}
   );
   gpc1_1 gpc1_1_4043(
      {stage127[111]},
      {stage127[195]}
   );
   gpc1_1 gpc1_1_4044(
      {stage127[112]},
      {stage127[196]}
   );
   gpc1_1 gpc1_1_4045(
      {stage127[113]},
      {stage127[197]}
   );
   gpc1_1 gpc1_1_4046(
      {stage127[114]},
      {stage127[198]}
   );
   gpc1_1 gpc1_1_4047(
      {stage127[115]},
      {stage127[199]}
   );
   gpc1_1 gpc1_1_4048(
      {stage127[116]},
      {stage127[200]}
   );
   gpc1_1 gpc1_1_4049(
      {stage127[117]},
      {stage127[201]}
   );
   gpc1_1 gpc1_1_4050(
      {stage127[118]},
      {stage127[202]}
   );
   gpc1_1 gpc1_1_4051(
      {stage127[119]},
      {stage127[203]}
   );
   gpc1_1 gpc1_1_4052(
      {stage127[120]},
      {stage127[204]}
   );
   gpc1_1 gpc1_1_4053(
      {stage127[121]},
      {stage127[205]}
   );
   gpc1_1 gpc1_1_4054(
      {stage127[122]},
      {stage127[206]}
   );
   gpc1_1 gpc1_1_4055(
      {stage127[123]},
      {stage127[207]}
   );
   gpc1_1 gpc1_1_4056(
      {stage127[124]},
      {stage127[208]}
   );
   gpc1_1 gpc1_1_4057(
      {stage127[125]},
      {stage127[209]}
   );
   gpc1_1 gpc1_1_4058(
      {stage127[126]},
      {stage127[210]}
   );
   gpc1_1 gpc1_1_4059(
      {stage127[127]},
      {stage127[211]}
   );
   gpc1_1 gpc1_1_4060(
      {stage000[128]},
      {stage000[170]}
   );
   gpc1_1 gpc1_1_4061(
      {stage000[129]},
      {stage000[171]}
   );
   gpc1_1 gpc1_1_4062(
      {stage000[130]},
      {stage000[172]}
   );
   gpc606_5 gpc606_5_4063(
      {stage000[131], stage000[132], stage000[133], stage000[134], stage000[135], stage000[136]},
      {stage002[128], stage002[129], stage002[130], stage002[131], stage002[132], stage002[133]},
      {stage004[186], stage003[176], stage002[189], stage001[183], stage000[173]}
   );
   gpc606_5 gpc606_5_4064(
      {stage000[137], stage000[138], stage000[139], stage000[140], stage000[141], stage000[142]},
      {stage002[134], stage002[135], stage002[136], stage002[137], stage002[138], stage002[139]},
      {stage004[187], stage003[177], stage002[190], stage001[184], stage000[174]}
   );
   gpc606_5 gpc606_5_4065(
      {stage000[143], stage000[144], stage000[145], stage000[146], stage000[147], stage000[148]},
      {stage002[140], stage002[141], stage002[142], stage002[143], stage002[144], stage002[145]},
      {stage004[188], stage003[178], stage002[191], stage001[185], stage000[175]}
   );
   gpc606_5 gpc606_5_4066(
      {stage000[149], stage000[150], stage000[151], stage000[152], stage000[153], stage000[154]},
      {stage002[146], stage002[147], stage002[148], stage002[149], stage002[150], stage002[151]},
      {stage004[189], stage003[179], stage002[192], stage001[186], stage000[176]}
   );
   gpc2135_5 gpc2135_5_4067(
      {stage000[155], stage000[156], stage000[157], stage000[158], stage000[159]},
      {stage001[128], stage001[129], stage001[130]},
      {stage002[152]},
      {stage003[128], stage003[129]},
      {stage004[190], stage003[180], stage002[193], stage001[187], stage000[177]}
   );
   gpc2135_5 gpc2135_5_4068(
      {stage000[160], stage000[161], stage000[162], stage000[163], stage000[164]},
      {stage001[131], stage001[132], stage001[133]},
      {stage002[153]},
      {stage003[130], stage003[131]},
      {stage004[191], stage003[181], stage002[194], stage001[188], stage000[178]}
   );
   gpc2135_5 gpc2135_5_4069(
      {stage000[165], stage000[166], stage000[167], stage000[168], stage000[169]},
      {stage001[134], stage001[135], stage001[136]},
      {stage002[154]},
      {stage003[132], stage003[133]},
      {stage004[192], stage003[182], stage002[195], stage001[189], stage000[179]}
   );
   gpc1_1 gpc1_1_4070(
      {stage001[137]},
      {stage001[190]}
   );
   gpc1_1 gpc1_1_4071(
      {stage001[138]},
      {stage001[191]}
   );
   gpc1_1 gpc1_1_4072(
      {stage001[139]},
      {stage001[192]}
   );
   gpc1_1 gpc1_1_4073(
      {stage001[140]},
      {stage001[193]}
   );
   gpc1_1 gpc1_1_4074(
      {stage001[141]},
      {stage001[194]}
   );
   gpc1_1 gpc1_1_4075(
      {stage001[142]},
      {stage001[195]}
   );
   gpc1_1 gpc1_1_4076(
      {stage001[143]},
      {stage001[196]}
   );
   gpc1_1 gpc1_1_4077(
      {stage001[144]},
      {stage001[197]}
   );
   gpc1_1 gpc1_1_4078(
      {stage001[145]},
      {stage001[198]}
   );
   gpc1_1 gpc1_1_4079(
      {stage001[146]},
      {stage001[199]}
   );
   gpc1_1 gpc1_1_4080(
      {stage001[147]},
      {stage001[200]}
   );
   gpc1_1 gpc1_1_4081(
      {stage001[148]},
      {stage001[201]}
   );
   gpc1_1 gpc1_1_4082(
      {stage001[149]},
      {stage001[202]}
   );
   gpc1_1 gpc1_1_4083(
      {stage001[150]},
      {stage001[203]}
   );
   gpc606_5 gpc606_5_4084(
      {stage001[151], stage001[152], stage001[153], stage001[154], stage001[155], stage001[156]},
      {stage003[134], stage003[135], stage003[136], stage003[137], stage003[138], stage003[139]},
      {stage005[213], stage004[193], stage003[183], stage002[196], stage001[204]}
   );
   gpc606_5 gpc606_5_4085(
      {stage001[157], stage001[158], stage001[159], stage001[160], stage001[161], stage001[162]},
      {stage003[140], stage003[141], stage003[142], stage003[143], stage003[144], stage003[145]},
      {stage005[214], stage004[194], stage003[184], stage002[197], stage001[205]}
   );
   gpc2135_5 gpc2135_5_4086(
      {stage001[163], stage001[164], stage001[165], stage001[166], stage001[167]},
      {stage002[155], stage002[156], stage002[157]},
      {stage003[146]},
      {stage004[128], stage004[129]},
      {stage005[215], stage004[195], stage003[185], stage002[198], stage001[206]}
   );
   gpc2135_5 gpc2135_5_4087(
      {stage001[168], stage001[169], stage001[170], stage001[171], stage001[172]},
      {stage002[158], stage002[159], stage002[160]},
      {stage003[147]},
      {stage004[130], stage004[131]},
      {stage005[216], stage004[196], stage003[186], stage002[199], stage001[207]}
   );
   gpc2135_5 gpc2135_5_4088(
      {stage001[173], stage001[174], stage001[175], stage001[176], stage001[177]},
      {stage002[161], stage002[162], stage002[163]},
      {stage003[148]},
      {stage004[132], stage004[133]},
      {stage005[217], stage004[197], stage003[187], stage002[200], stage001[208]}
   );
   gpc2135_5 gpc2135_5_4089(
      {stage001[178], stage001[179], stage001[180], stage001[181], stage001[182]},
      {stage002[164], stage002[165], stage002[166]},
      {stage003[149]},
      {stage004[134], stage004[135]},
      {stage005[218], stage004[198], stage003[188], stage002[201], stage001[209]}
   );
   gpc1_1 gpc1_1_4090(
      {stage002[167]},
      {stage002[202]}
   );
   gpc1_1 gpc1_1_4091(
      {stage002[168]},
      {stage002[203]}
   );
   gpc1_1 gpc1_1_4092(
      {stage002[169]},
      {stage002[204]}
   );
   gpc1_1 gpc1_1_4093(
      {stage002[170]},
      {stage002[205]}
   );
   gpc1_1 gpc1_1_4094(
      {stage002[171]},
      {stage002[206]}
   );
   gpc1_1 gpc1_1_4095(
      {stage002[172]},
      {stage002[207]}
   );
   gpc1_1 gpc1_1_4096(
      {stage002[173]},
      {stage002[208]}
   );
   gpc1_1 gpc1_1_4097(
      {stage002[174]},
      {stage002[209]}
   );
   gpc1_1 gpc1_1_4098(
      {stage002[175]},
      {stage002[210]}
   );
   gpc1_1 gpc1_1_4099(
      {stage002[176]},
      {stage002[211]}
   );
   gpc1_1 gpc1_1_4100(
      {stage002[177]},
      {stage002[212]}
   );
   gpc1_1 gpc1_1_4101(
      {stage002[178]},
      {stage002[213]}
   );
   gpc1_1 gpc1_1_4102(
      {stage002[179]},
      {stage002[214]}
   );
   gpc1_1 gpc1_1_4103(
      {stage002[180]},
      {stage002[215]}
   );
   gpc1_1 gpc1_1_4104(
      {stage002[181]},
      {stage002[216]}
   );
   gpc1_1 gpc1_1_4105(
      {stage002[182]},
      {stage002[217]}
   );
   gpc606_5 gpc606_5_4106(
      {stage002[183], stage002[184], stage002[185], stage002[186], stage002[187], stage002[188]},
      {stage004[136], stage004[137], stage004[138], stage004[139], stage004[140], stage004[141]},
      {stage006[188], stage005[219], stage004[199], stage003[189], stage002[218]}
   );
   gpc623_5 gpc623_5_4107(
      {stage003[150], stage003[151], stage003[152]},
      {stage004[142], stage004[143]},
      {stage005[128], stage005[129], stage005[130], stage005[131], stage005[132], stage005[133]},
      {stage007[193], stage006[189], stage005[220], stage004[200], stage003[190]}
   );
   gpc623_5 gpc623_5_4108(
      {stage003[153], stage003[154], stage003[155]},
      {stage004[144], stage004[145]},
      {stage005[134], stage005[135], stage005[136], stage005[137], stage005[138], stage005[139]},
      {stage007[194], stage006[190], stage005[221], stage004[201], stage003[191]}
   );
   gpc623_5 gpc623_5_4109(
      {stage003[156], stage003[157], stage003[158]},
      {stage004[146], stage004[147]},
      {stage005[140], stage005[141], stage005[142], stage005[143], stage005[144], stage005[145]},
      {stage007[195], stage006[191], stage005[222], stage004[202], stage003[192]}
   );
   gpc623_5 gpc623_5_4110(
      {stage003[159], stage003[160], stage003[161]},
      {stage004[148], stage004[149]},
      {stage005[146], stage005[147], stage005[148], stage005[149], stage005[150], stage005[151]},
      {stage007[196], stage006[192], stage005[223], stage004[203], stage003[193]}
   );
   gpc615_5 gpc615_5_4111(
      {stage003[162], stage003[163], stage003[164], stage003[165], stage003[166]},
      {stage004[150]},
      {stage005[152], stage005[153], stage005[154], stage005[155], stage005[156], stage005[157]},
      {stage007[197], stage006[193], stage005[224], stage004[204], stage003[194]}
   );
   gpc615_5 gpc615_5_4112(
      {stage003[167], stage003[168], stage003[169], stage003[170], stage003[171]},
      {stage004[151]},
      {stage005[158], stage005[159], stage005[160], stage005[161], stage005[162], stage005[163]},
      {stage007[198], stage006[194], stage005[225], stage004[205], stage003[195]}
   );
   gpc615_5 gpc615_5_4113(
      {stage003[172], stage003[173], stage003[174], stage003[175], 1'h0},
      {stage004[152]},
      {stage005[164], stage005[165], stage005[166], stage005[167], stage005[168], stage005[169]},
      {stage007[199], stage006[195], stage005[226], stage004[206], stage003[196]}
   );
   gpc1_1 gpc1_1_4114(
      {stage004[153]},
      {stage004[207]}
   );
   gpc1_1 gpc1_1_4115(
      {stage004[154]},
      {stage004[208]}
   );
   gpc1_1 gpc1_1_4116(
      {stage004[155]},
      {stage004[209]}
   );
   gpc1_1 gpc1_1_4117(
      {stage004[156]},
      {stage004[210]}
   );
   gpc1_1 gpc1_1_4118(
      {stage004[157]},
      {stage004[211]}
   );
   gpc1_1 gpc1_1_4119(
      {stage004[158]},
      {stage004[212]}
   );
   gpc1_1 gpc1_1_4120(
      {stage004[159]},
      {stage004[213]}
   );
   gpc1_1 gpc1_1_4121(
      {stage004[160]},
      {stage004[214]}
   );
   gpc1_1 gpc1_1_4122(
      {stage004[161]},
      {stage004[215]}
   );
   gpc1_1 gpc1_1_4123(
      {stage004[162]},
      {stage004[216]}
   );
   gpc1_1 gpc1_1_4124(
      {stage004[163]},
      {stage004[217]}
   );
   gpc1_1 gpc1_1_4125(
      {stage004[164]},
      {stage004[218]}
   );
   gpc1_1 gpc1_1_4126(
      {stage004[165]},
      {stage004[219]}
   );
   gpc1_1 gpc1_1_4127(
      {stage004[166]},
      {stage004[220]}
   );
   gpc1_1 gpc1_1_4128(
      {stage004[167]},
      {stage004[221]}
   );
   gpc1_1 gpc1_1_4129(
      {stage004[168]},
      {stage004[222]}
   );
   gpc1_1 gpc1_1_4130(
      {stage004[169]},
      {stage004[223]}
   );
   gpc1_1 gpc1_1_4131(
      {stage004[170]},
      {stage004[224]}
   );
   gpc1_1 gpc1_1_4132(
      {stage004[171]},
      {stage004[225]}
   );
   gpc1_1 gpc1_1_4133(
      {stage004[172]},
      {stage004[226]}
   );
   gpc1_1 gpc1_1_4134(
      {stage004[173]},
      {stage004[227]}
   );
   gpc1_1 gpc1_1_4135(
      {stage004[174]},
      {stage004[228]}
   );
   gpc1_1 gpc1_1_4136(
      {stage004[175]},
      {stage004[229]}
   );
   gpc615_5 gpc615_5_4137(
      {stage004[176], stage004[177], stage004[178], stage004[179], stage004[180]},
      {stage005[170]},
      {stage006[128], stage006[129], stage006[130], stage006[131], stage006[132], stage006[133]},
      {stage008[176], stage007[200], stage006[196], stage005[227], stage004[230]}
   );
   gpc615_5 gpc615_5_4138(
      {stage004[181], stage004[182], stage004[183], stage004[184], stage004[185]},
      {stage005[171]},
      {stage006[134], stage006[135], stage006[136], stage006[137], stage006[138], stage006[139]},
      {stage008[177], stage007[201], stage006[197], stage005[228], stage004[231]}
   );
   gpc1_1 gpc1_1_4139(
      {stage005[172]},
      {stage005[229]}
   );
   gpc1_1 gpc1_1_4140(
      {stage005[173]},
      {stage005[230]}
   );
   gpc1_1 gpc1_1_4141(
      {stage005[174]},
      {stage005[231]}
   );
   gpc1_1 gpc1_1_4142(
      {stage005[175]},
      {stage005[232]}
   );
   gpc1_1 gpc1_1_4143(
      {stage005[176]},
      {stage005[233]}
   );
   gpc1_1 gpc1_1_4144(
      {stage005[177]},
      {stage005[234]}
   );
   gpc1_1 gpc1_1_4145(
      {stage005[178]},
      {stage005[235]}
   );
   gpc1_1 gpc1_1_4146(
      {stage005[179]},
      {stage005[236]}
   );
   gpc1_1 gpc1_1_4147(
      {stage005[180]},
      {stage005[237]}
   );
   gpc1_1 gpc1_1_4148(
      {stage005[181]},
      {stage005[238]}
   );
   gpc1_1 gpc1_1_4149(
      {stage005[182]},
      {stage005[239]}
   );
   gpc606_5 gpc606_5_4150(
      {stage005[183], stage005[184], stage005[185], stage005[186], stage005[187], stage005[188]},
      {stage007[128], stage007[129], stage007[130], stage007[131], stage007[132], stage007[133]},
      {stage009[188], stage008[178], stage007[202], stage006[198], stage005[240]}
   );
   gpc606_5 gpc606_5_4151(
      {stage005[189], stage005[190], stage005[191], stage005[192], stage005[193], stage005[194]},
      {stage007[134], stage007[135], stage007[136], stage007[137], stage007[138], stage007[139]},
      {stage009[189], stage008[179], stage007[203], stage006[199], stage005[241]}
   );
   gpc606_5 gpc606_5_4152(
      {stage005[195], stage005[196], stage005[197], stage005[198], stage005[199], stage005[200]},
      {stage007[140], stage007[141], stage007[142], stage007[143], stage007[144], stage007[145]},
      {stage009[190], stage008[180], stage007[204], stage006[200], stage005[242]}
   );
   gpc606_5 gpc606_5_4153(
      {stage005[201], stage005[202], stage005[203], stage005[204], stage005[205], stage005[206]},
      {stage007[146], stage007[147], stage007[148], stage007[149], stage007[150], stage007[151]},
      {stage009[191], stage008[181], stage007[205], stage006[201], stage005[243]}
   );
   gpc606_5 gpc606_5_4154(
      {stage005[207], stage005[208], stage005[209], stage005[210], stage005[211], stage005[212]},
      {stage007[152], stage007[153], stage007[154], stage007[155], stage007[156], stage007[157]},
      {stage009[192], stage008[182], stage007[206], stage006[202], stage005[244]}
   );
   gpc1_1 gpc1_1_4155(
      {stage006[140]},
      {stage006[203]}
   );
   gpc1_1 gpc1_1_4156(
      {stage006[141]},
      {stage006[204]}
   );
   gpc1_1 gpc1_1_4157(
      {stage006[142]},
      {stage006[205]}
   );
   gpc1_1 gpc1_1_4158(
      {stage006[143]},
      {stage006[206]}
   );
   gpc1_1 gpc1_1_4159(
      {stage006[144]},
      {stage006[207]}
   );
   gpc1_1 gpc1_1_4160(
      {stage006[145]},
      {stage006[208]}
   );
   gpc1_1 gpc1_1_4161(
      {stage006[146]},
      {stage006[209]}
   );
   gpc1_1 gpc1_1_4162(
      {stage006[147]},
      {stage006[210]}
   );
   gpc1_1 gpc1_1_4163(
      {stage006[148]},
      {stage006[211]}
   );
   gpc1_1 gpc1_1_4164(
      {stage006[149]},
      {stage006[212]}
   );
   gpc1_1 gpc1_1_4165(
      {stage006[150]},
      {stage006[213]}
   );
   gpc1_1 gpc1_1_4166(
      {stage006[151]},
      {stage006[214]}
   );
   gpc1_1 gpc1_1_4167(
      {stage006[152]},
      {stage006[215]}
   );
   gpc1_1 gpc1_1_4168(
      {stage006[153]},
      {stage006[216]}
   );
   gpc1_1 gpc1_1_4169(
      {stage006[154]},
      {stage006[217]}
   );
   gpc1_1 gpc1_1_4170(
      {stage006[155]},
      {stage006[218]}
   );
   gpc1_1 gpc1_1_4171(
      {stage006[156]},
      {stage006[219]}
   );
   gpc1_1 gpc1_1_4172(
      {stage006[157]},
      {stage006[220]}
   );
   gpc606_5 gpc606_5_4173(
      {stage006[158], stage006[159], stage006[160], stage006[161], stage006[162], stage006[163]},
      {stage008[128], stage008[129], stage008[130], stage008[131], stage008[132], stage008[133]},
      {stage010[188], stage009[193], stage008[183], stage007[207], stage006[221]}
   );
   gpc606_5 gpc606_5_4174(
      {stage006[164], stage006[165], stage006[166], stage006[167], stage006[168], stage006[169]},
      {stage008[134], stage008[135], stage008[136], stage008[137], stage008[138], stage008[139]},
      {stage010[189], stage009[194], stage008[184], stage007[208], stage006[222]}
   );
   gpc606_5 gpc606_5_4175(
      {stage006[170], stage006[171], stage006[172], stage006[173], stage006[174], stage006[175]},
      {stage008[140], stage008[141], stage008[142], stage008[143], stage008[144], stage008[145]},
      {stage010[190], stage009[195], stage008[185], stage007[209], stage006[223]}
   );
   gpc606_5 gpc606_5_4176(
      {stage006[176], stage006[177], stage006[178], stage006[179], stage006[180], stage006[181]},
      {stage008[146], stage008[147], stage008[148], stage008[149], stage008[150], stage008[151]},
      {stage010[191], stage009[196], stage008[186], stage007[210], stage006[224]}
   );
   gpc606_5 gpc606_5_4177(
      {stage006[182], stage006[183], stage006[184], stage006[185], stage006[186], stage006[187]},
      {stage008[152], stage008[153], stage008[154], stage008[155], stage008[156], stage008[157]},
      {stage010[192], stage009[197], stage008[187], stage007[211], stage006[225]}
   );
   gpc1_1 gpc1_1_4178(
      {stage007[158]},
      {stage007[212]}
   );
   gpc1_1 gpc1_1_4179(
      {stage007[159]},
      {stage007[213]}
   );
   gpc1_1 gpc1_1_4180(
      {stage007[160]},
      {stage007[214]}
   );
   gpc1_1 gpc1_1_4181(
      {stage007[161]},
      {stage007[215]}
   );
   gpc1_1 gpc1_1_4182(
      {stage007[162]},
      {stage007[216]}
   );
   gpc1_1 gpc1_1_4183(
      {stage007[163]},
      {stage007[217]}
   );
   gpc1_1 gpc1_1_4184(
      {stage007[164]},
      {stage007[218]}
   );
   gpc1_1 gpc1_1_4185(
      {stage007[165]},
      {stage007[219]}
   );
   gpc1_1 gpc1_1_4186(
      {stage007[166]},
      {stage007[220]}
   );
   gpc1_1 gpc1_1_4187(
      {stage007[167]},
      {stage007[221]}
   );
   gpc1_1 gpc1_1_4188(
      {stage007[168]},
      {stage007[222]}
   );
   gpc1_1 gpc1_1_4189(
      {stage007[169]},
      {stage007[223]}
   );
   gpc606_5 gpc606_5_4190(
      {stage007[170], stage007[171], stage007[172], stage007[173], stage007[174], stage007[175]},
      {stage009[128], stage009[129], stage009[130], stage009[131], stage009[132], stage009[133]},
      {stage011[202], stage010[193], stage009[198], stage008[188], stage007[224]}
   );
   gpc606_5 gpc606_5_4191(
      {stage007[176], stage007[177], stage007[178], stage007[179], stage007[180], stage007[181]},
      {stage009[134], stage009[135], stage009[136], stage009[137], stage009[138], stage009[139]},
      {stage011[203], stage010[194], stage009[199], stage008[189], stage007[225]}
   );
   gpc606_5 gpc606_5_4192(
      {stage007[182], stage007[183], stage007[184], stage007[185], stage007[186], stage007[187]},
      {stage009[140], stage009[141], stage009[142], stage009[143], stage009[144], stage009[145]},
      {stage011[204], stage010[195], stage009[200], stage008[190], stage007[226]}
   );
   gpc615_5 gpc615_5_4193(
      {stage007[188], stage007[189], stage007[190], stage007[191], stage007[192]},
      {stage008[158]},
      {stage009[146], stage009[147], stage009[148], stage009[149], stage009[150], stage009[151]},
      {stage011[205], stage010[196], stage009[201], stage008[191], stage007[227]}
   );
   gpc1_1 gpc1_1_4194(
      {stage008[159]},
      {stage008[192]}
   );
   gpc1_1 gpc1_1_4195(
      {stage008[160]},
      {stage008[193]}
   );
   gpc1_1 gpc1_1_4196(
      {stage008[161]},
      {stage008[194]}
   );
   gpc1_1 gpc1_1_4197(
      {stage008[162]},
      {stage008[195]}
   );
   gpc1_1 gpc1_1_4198(
      {stage008[163]},
      {stage008[196]}
   );
   gpc1_1 gpc1_1_4199(
      {stage008[164]},
      {stage008[197]}
   );
   gpc1_1 gpc1_1_4200(
      {stage008[165]},
      {stage008[198]}
   );
   gpc1_1 gpc1_1_4201(
      {stage008[166]},
      {stage008[199]}
   );
   gpc1_1 gpc1_1_4202(
      {stage008[167]},
      {stage008[200]}
   );
   gpc1_1 gpc1_1_4203(
      {stage008[168]},
      {stage008[201]}
   );
   gpc1_1 gpc1_1_4204(
      {stage008[169]},
      {stage008[202]}
   );
   gpc1_1 gpc1_1_4205(
      {stage008[170]},
      {stage008[203]}
   );
   gpc615_5 gpc615_5_4206(
      {stage008[171], stage008[172], stage008[173], stage008[174], stage008[175]},
      {stage009[152]},
      {stage010[128], stage010[129], stage010[130], stage010[131], stage010[132], stage010[133]},
      {stage012[220], stage011[206], stage010[197], stage009[202], stage008[204]}
   );
   gpc1_1 gpc1_1_4207(
      {stage009[153]},
      {stage009[203]}
   );
   gpc1_1 gpc1_1_4208(
      {stage009[154]},
      {stage009[204]}
   );
   gpc1_1 gpc1_1_4209(
      {stage009[155]},
      {stage009[205]}
   );
   gpc1_1 gpc1_1_4210(
      {stage009[156]},
      {stage009[206]}
   );
   gpc1_1 gpc1_1_4211(
      {stage009[157]},
      {stage009[207]}
   );
   gpc606_5 gpc606_5_4212(
      {stage009[158], stage009[159], stage009[160], stage009[161], stage009[162], stage009[163]},
      {stage011[128], stage011[129], stage011[130], stage011[131], stage011[132], stage011[133]},
      {stage013[184], stage012[221], stage011[207], stage010[198], stage009[208]}
   );
   gpc606_5 gpc606_5_4213(
      {stage009[164], stage009[165], stage009[166], stage009[167], stage009[168], stage009[169]},
      {stage011[134], stage011[135], stage011[136], stage011[137], stage011[138], stage011[139]},
      {stage013[185], stage012[222], stage011[208], stage010[199], stage009[209]}
   );
   gpc606_5 gpc606_5_4214(
      {stage009[170], stage009[171], stage009[172], stage009[173], stage009[174], stage009[175]},
      {stage011[140], stage011[141], stage011[142], stage011[143], stage011[144], stage011[145]},
      {stage013[186], stage012[223], stage011[209], stage010[200], stage009[210]}
   );
   gpc606_5 gpc606_5_4215(
      {stage009[176], stage009[177], stage009[178], stage009[179], stage009[180], stage009[181]},
      {stage011[146], stage011[147], stage011[148], stage011[149], stage011[150], stage011[151]},
      {stage013[187], stage012[224], stage011[210], stage010[201], stage009[211]}
   );
   gpc606_5 gpc606_5_4216(
      {stage009[182], stage009[183], stage009[184], stage009[185], stage009[186], stage009[187]},
      {stage011[152], stage011[153], stage011[154], stage011[155], stage011[156], stage011[157]},
      {stage013[188], stage012[225], stage011[211], stage010[202], stage009[212]}
   );
   gpc1_1 gpc1_1_4217(
      {stage010[134]},
      {stage010[203]}
   );
   gpc1_1 gpc1_1_4218(
      {stage010[135]},
      {stage010[204]}
   );
   gpc1_1 gpc1_1_4219(
      {stage010[136]},
      {stage010[205]}
   );
   gpc1_1 gpc1_1_4220(
      {stage010[137]},
      {stage010[206]}
   );
   gpc1_1 gpc1_1_4221(
      {stage010[138]},
      {stage010[207]}
   );
   gpc1_1 gpc1_1_4222(
      {stage010[139]},
      {stage010[208]}
   );
   gpc1_1 gpc1_1_4223(
      {stage010[140]},
      {stage010[209]}
   );
   gpc1_1 gpc1_1_4224(
      {stage010[141]},
      {stage010[210]}
   );
   gpc1_1 gpc1_1_4225(
      {stage010[142]},
      {stage010[211]}
   );
   gpc1_1 gpc1_1_4226(
      {stage010[143]},
      {stage010[212]}
   );
   gpc1_1 gpc1_1_4227(
      {stage010[144]},
      {stage010[213]}
   );
   gpc1_1 gpc1_1_4228(
      {stage010[145]},
      {stage010[214]}
   );
   gpc1_1 gpc1_1_4229(
      {stage010[146]},
      {stage010[215]}
   );
   gpc1_1 gpc1_1_4230(
      {stage010[147]},
      {stage010[216]}
   );
   gpc1_1 gpc1_1_4231(
      {stage010[148]},
      {stage010[217]}
   );
   gpc1_1 gpc1_1_4232(
      {stage010[149]},
      {stage010[218]}
   );
   gpc1_1 gpc1_1_4233(
      {stage010[150]},
      {stage010[219]}
   );
   gpc1_1 gpc1_1_4234(
      {stage010[151]},
      {stage010[220]}
   );
   gpc1_1 gpc1_1_4235(
      {stage010[152]},
      {stage010[221]}
   );
   gpc1_1 gpc1_1_4236(
      {stage010[153]},
      {stage010[222]}
   );
   gpc1_1 gpc1_1_4237(
      {stage010[154]},
      {stage010[223]}
   );
   gpc1_1 gpc1_1_4238(
      {stage010[155]},
      {stage010[224]}
   );
   gpc1_1 gpc1_1_4239(
      {stage010[156]},
      {stage010[225]}
   );
   gpc1_1 gpc1_1_4240(
      {stage010[157]},
      {stage010[226]}
   );
   gpc1_1 gpc1_1_4241(
      {stage010[158]},
      {stage010[227]}
   );
   gpc1_1 gpc1_1_4242(
      {stage010[159]},
      {stage010[228]}
   );
   gpc1_1 gpc1_1_4243(
      {stage010[160]},
      {stage010[229]}
   );
   gpc1_1 gpc1_1_4244(
      {stage010[161]},
      {stage010[230]}
   );
   gpc1_1 gpc1_1_4245(
      {stage010[162]},
      {stage010[231]}
   );
   gpc1_1 gpc1_1_4246(
      {stage010[163]},
      {stage010[232]}
   );
   gpc1_1 gpc1_1_4247(
      {stage010[164]},
      {stage010[233]}
   );
   gpc1_1 gpc1_1_4248(
      {stage010[165]},
      {stage010[234]}
   );
   gpc1_1 gpc1_1_4249(
      {stage010[166]},
      {stage010[235]}
   );
   gpc1_1 gpc1_1_4250(
      {stage010[167]},
      {stage010[236]}
   );
   gpc1_1 gpc1_1_4251(
      {stage010[168]},
      {stage010[237]}
   );
   gpc1_1 gpc1_1_4252(
      {stage010[169]},
      {stage010[238]}
   );
   gpc1_1 gpc1_1_4253(
      {stage010[170]},
      {stage010[239]}
   );
   gpc1_1 gpc1_1_4254(
      {stage010[171]},
      {stage010[240]}
   );
   gpc1_1 gpc1_1_4255(
      {stage010[172]},
      {stage010[241]}
   );
   gpc1_1 gpc1_1_4256(
      {stage010[173]},
      {stage010[242]}
   );
   gpc1_1 gpc1_1_4257(
      {stage010[174]},
      {stage010[243]}
   );
   gpc1_1 gpc1_1_4258(
      {stage010[175]},
      {stage010[244]}
   );
   gpc1_1 gpc1_1_4259(
      {stage010[176]},
      {stage010[245]}
   );
   gpc1_1 gpc1_1_4260(
      {stage010[177]},
      {stage010[246]}
   );
   gpc1_1 gpc1_1_4261(
      {stage010[178]},
      {stage010[247]}
   );
   gpc1_1 gpc1_1_4262(
      {stage010[179]},
      {stage010[248]}
   );
   gpc1_1 gpc1_1_4263(
      {stage010[180]},
      {stage010[249]}
   );
   gpc1_1 gpc1_1_4264(
      {stage010[181]},
      {stage010[250]}
   );
   gpc1_1 gpc1_1_4265(
      {stage010[182]},
      {stage010[251]}
   );
   gpc1_1 gpc1_1_4266(
      {stage010[183]},
      {stage010[252]}
   );
   gpc1_1 gpc1_1_4267(
      {stage010[184]},
      {stage010[253]}
   );
   gpc1_1 gpc1_1_4268(
      {stage010[185]},
      {stage010[254]}
   );
   gpc1_1 gpc1_1_4269(
      {stage010[186]},
      {stage010[255]}
   );
   gpc1_1 gpc1_1_4270(
      {stage010[187]},
      {stage010[256]}
   );
   gpc606_5 gpc606_5_4271(
      {stage011[158], stage011[159], stage011[160], stage011[161], stage011[162], stage011[163]},
      {stage013[128], stage013[129], stage013[130], stage013[131], stage013[132], stage013[133]},
      {stage015[188], stage014[227], stage013[189], stage012[226], stage011[212]}
   );
   gpc606_5 gpc606_5_4272(
      {stage011[164], stage011[165], stage011[166], stage011[167], stage011[168], stage011[169]},
      {stage013[134], stage013[135], stage013[136], stage013[137], stage013[138], stage013[139]},
      {stage015[189], stage014[228], stage013[190], stage012[227], stage011[213]}
   );
   gpc606_5 gpc606_5_4273(
      {stage011[170], stage011[171], stage011[172], stage011[173], stage011[174], stage011[175]},
      {stage013[140], stage013[141], stage013[142], stage013[143], stage013[144], stage013[145]},
      {stage015[190], stage014[229], stage013[191], stage012[228], stage011[214]}
   );
   gpc606_5 gpc606_5_4274(
      {stage011[176], stage011[177], stage011[178], stage011[179], stage011[180], stage011[181]},
      {stage013[146], stage013[147], stage013[148], stage013[149], stage013[150], stage013[151]},
      {stage015[191], stage014[230], stage013[192], stage012[229], stage011[215]}
   );
   gpc615_5 gpc615_5_4275(
      {stage011[182], stage011[183], stage011[184], stage011[185], stage011[186]},
      {stage012[128]},
      {stage013[152], stage013[153], stage013[154], stage013[155], stage013[156], stage013[157]},
      {stage015[192], stage014[231], stage013[193], stage012[230], stage011[216]}
   );
   gpc615_5 gpc615_5_4276(
      {stage011[187], stage011[188], stage011[189], stage011[190], stage011[191]},
      {stage012[129]},
      {stage013[158], stage013[159], stage013[160], stage013[161], stage013[162], stage013[163]},
      {stage015[193], stage014[232], stage013[194], stage012[231], stage011[217]}
   );
   gpc615_5 gpc615_5_4277(
      {stage011[192], stage011[193], stage011[194], stage011[195], stage011[196]},
      {stage012[130]},
      {stage013[164], stage013[165], stage013[166], stage013[167], stage013[168], stage013[169]},
      {stage015[194], stage014[233], stage013[195], stage012[232], stage011[218]}
   );
   gpc1325_5 gpc1325_5_4278(
      {stage011[197], stage011[198], stage011[199], stage011[200], stage011[201]},
      {stage012[131], stage012[132]},
      {stage013[170], stage013[171], stage013[172]},
      {stage014[128]},
      {stage015[195], stage014[234], stage013[196], stage012[233], stage011[219]}
   );
   gpc1_1 gpc1_1_4279(
      {stage012[133]},
      {stage012[234]}
   );
   gpc1_1 gpc1_1_4280(
      {stage012[134]},
      {stage012[235]}
   );
   gpc1_1 gpc1_1_4281(
      {stage012[135]},
      {stage012[236]}
   );
   gpc1_1 gpc1_1_4282(
      {stage012[136]},
      {stage012[237]}
   );
   gpc1_1 gpc1_1_4283(
      {stage012[137]},
      {stage012[238]}
   );
   gpc1_1 gpc1_1_4284(
      {stage012[138]},
      {stage012[239]}
   );
   gpc1_1 gpc1_1_4285(
      {stage012[139]},
      {stage012[240]}
   );
   gpc1_1 gpc1_1_4286(
      {stage012[140]},
      {stage012[241]}
   );
   gpc1_1 gpc1_1_4287(
      {stage012[141]},
      {stage012[242]}
   );
   gpc1_1 gpc1_1_4288(
      {stage012[142]},
      {stage012[243]}
   );
   gpc1_1 gpc1_1_4289(
      {stage012[143]},
      {stage012[244]}
   );
   gpc1_1 gpc1_1_4290(
      {stage012[144]},
      {stage012[245]}
   );
   gpc1_1 gpc1_1_4291(
      {stage012[145]},
      {stage012[246]}
   );
   gpc1_1 gpc1_1_4292(
      {stage012[146]},
      {stage012[247]}
   );
   gpc1_1 gpc1_1_4293(
      {stage012[147]},
      {stage012[248]}
   );
   gpc1_1 gpc1_1_4294(
      {stage012[148]},
      {stage012[249]}
   );
   gpc1_1 gpc1_1_4295(
      {stage012[149]},
      {stage012[250]}
   );
   gpc1_1 gpc1_1_4296(
      {stage012[150]},
      {stage012[251]}
   );
   gpc1_1 gpc1_1_4297(
      {stage012[151]},
      {stage012[252]}
   );
   gpc1_1 gpc1_1_4298(
      {stage012[152]},
      {stage012[253]}
   );
   gpc1_1 gpc1_1_4299(
      {stage012[153]},
      {stage012[254]}
   );
   gpc1_1 gpc1_1_4300(
      {stage012[154]},
      {stage012[255]}
   );
   gpc1_1 gpc1_1_4301(
      {stage012[155]},
      {stage012[256]}
   );
   gpc1_1 gpc1_1_4302(
      {stage012[156]},
      {stage012[257]}
   );
   gpc1_1 gpc1_1_4303(
      {stage012[157]},
      {stage012[258]}
   );
   gpc1_1 gpc1_1_4304(
      {stage012[158]},
      {stage012[259]}
   );
   gpc1_1 gpc1_1_4305(
      {stage012[159]},
      {stage012[260]}
   );
   gpc1_1 gpc1_1_4306(
      {stage012[160]},
      {stage012[261]}
   );
   gpc1_1 gpc1_1_4307(
      {stage012[161]},
      {stage012[262]}
   );
   gpc1_1 gpc1_1_4308(
      {stage012[162]},
      {stage012[263]}
   );
   gpc1_1 gpc1_1_4309(
      {stage012[163]},
      {stage012[264]}
   );
   gpc1_1 gpc1_1_4310(
      {stage012[164]},
      {stage012[265]}
   );
   gpc615_5 gpc615_5_4311(
      {stage012[165], stage012[166], stage012[167], stage012[168], stage012[169]},
      {stage013[173]},
      {stage014[129], stage014[130], stage014[131], stage014[132], stage014[133], stage014[134]},
      {stage016[209], stage015[196], stage014[235], stage013[197], stage012[266]}
   );
   gpc615_5 gpc615_5_4312(
      {stage012[170], stage012[171], stage012[172], stage012[173], stage012[174]},
      {stage013[174]},
      {stage014[135], stage014[136], stage014[137], stage014[138], stage014[139], stage014[140]},
      {stage016[210], stage015[197], stage014[236], stage013[198], stage012[267]}
   );
   gpc615_5 gpc615_5_4313(
      {stage012[175], stage012[176], stage012[177], stage012[178], stage012[179]},
      {stage013[175]},
      {stage014[141], stage014[142], stage014[143], stage014[144], stage014[145], stage014[146]},
      {stage016[211], stage015[198], stage014[237], stage013[199], stage012[268]}
   );
   gpc615_5 gpc615_5_4314(
      {stage012[180], stage012[181], stage012[182], stage012[183], stage012[184]},
      {stage013[176]},
      {stage014[147], stage014[148], stage014[149], stage014[150], stage014[151], stage014[152]},
      {stage016[212], stage015[199], stage014[238], stage013[200], stage012[269]}
   );
   gpc615_5 gpc615_5_4315(
      {stage012[185], stage012[186], stage012[187], stage012[188], stage012[189]},
      {stage013[177]},
      {stage014[153], stage014[154], stage014[155], stage014[156], stage014[157], stage014[158]},
      {stage016[213], stage015[200], stage014[239], stage013[201], stage012[270]}
   );
   gpc615_5 gpc615_5_4316(
      {stage012[190], stage012[191], stage012[192], stage012[193], stage012[194]},
      {stage013[178]},
      {stage014[159], stage014[160], stage014[161], stage014[162], stage014[163], stage014[164]},
      {stage016[214], stage015[201], stage014[240], stage013[202], stage012[271]}
   );
   gpc615_5 gpc615_5_4317(
      {stage012[195], stage012[196], stage012[197], stage012[198], stage012[199]},
      {stage013[179]},
      {stage014[165], stage014[166], stage014[167], stage014[168], stage014[169], stage014[170]},
      {stage016[215], stage015[202], stage014[241], stage013[203], stage012[272]}
   );
   gpc615_5 gpc615_5_4318(
      {stage012[200], stage012[201], stage012[202], stage012[203], stage012[204]},
      {stage013[180]},
      {stage014[171], stage014[172], stage014[173], stage014[174], stage014[175], stage014[176]},
      {stage016[216], stage015[203], stage014[242], stage013[204], stage012[273]}
   );
   gpc615_5 gpc615_5_4319(
      {stage012[205], stage012[206], stage012[207], stage012[208], stage012[209]},
      {stage013[181]},
      {stage014[177], stage014[178], stage014[179], stage014[180], stage014[181], stage014[182]},
      {stage016[217], stage015[204], stage014[243], stage013[205], stage012[274]}
   );
   gpc615_5 gpc615_5_4320(
      {stage012[210], stage012[211], stage012[212], stage012[213], stage012[214]},
      {stage013[182]},
      {stage014[183], stage014[184], stage014[185], stage014[186], stage014[187], stage014[188]},
      {stage016[218], stage015[205], stage014[244], stage013[206], stage012[275]}
   );
   gpc615_5 gpc615_5_4321(
      {stage012[215], stage012[216], stage012[217], stage012[218], stage012[219]},
      {stage013[183]},
      {stage014[189], stage014[190], stage014[191], stage014[192], stage014[193], stage014[194]},
      {stage016[219], stage015[206], stage014[245], stage013[207], stage012[276]}
   );
   gpc1_1 gpc1_1_4322(
      {stage014[195]},
      {stage014[246]}
   );
   gpc1_1 gpc1_1_4323(
      {stage014[196]},
      {stage014[247]}
   );
   gpc1_1 gpc1_1_4324(
      {stage014[197]},
      {stage014[248]}
   );
   gpc1_1 gpc1_1_4325(
      {stage014[198]},
      {stage014[249]}
   );
   gpc1_1 gpc1_1_4326(
      {stage014[199]},
      {stage014[250]}
   );
   gpc1_1 gpc1_1_4327(
      {stage014[200]},
      {stage014[251]}
   );
   gpc1_1 gpc1_1_4328(
      {stage014[201]},
      {stage014[252]}
   );
   gpc1_1 gpc1_1_4329(
      {stage014[202]},
      {stage014[253]}
   );
   gpc606_5 gpc606_5_4330(
      {stage014[203], stage014[204], stage014[205], stage014[206], stage014[207], stage014[208]},
      {stage016[128], stage016[129], stage016[130], stage016[131], stage016[132], stage016[133]},
      {stage018[189], stage017[219], stage016[220], stage015[207], stage014[254]}
   );
   gpc606_5 gpc606_5_4331(
      {stage014[209], stage014[210], stage014[211], stage014[212], stage014[213], stage014[214]},
      {stage016[134], stage016[135], stage016[136], stage016[137], stage016[138], stage016[139]},
      {stage018[190], stage017[220], stage016[221], stage015[208], stage014[255]}
   );
   gpc606_5 gpc606_5_4332(
      {stage014[215], stage014[216], stage014[217], stage014[218], stage014[219], stage014[220]},
      {stage016[140], stage016[141], stage016[142], stage016[143], stage016[144], stage016[145]},
      {stage018[191], stage017[221], stage016[222], stage015[209], stage014[256]}
   );
   gpc606_5 gpc606_5_4333(
      {stage014[221], stage014[222], stage014[223], stage014[224], stage014[225], stage014[226]},
      {stage016[146], stage016[147], stage016[148], stage016[149], stage016[150], stage016[151]},
      {stage018[192], stage017[222], stage016[223], stage015[210], stage014[257]}
   );
   gpc615_5 gpc615_5_4334(
      {stage015[128], stage015[129], stage015[130], stage015[131], stage015[132]},
      {stage016[152]},
      {stage017[128], stage017[129], stage017[130], stage017[131], stage017[132], stage017[133]},
      {stage019[188], stage018[193], stage017[223], stage016[224], stage015[211]}
   );
   gpc615_5 gpc615_5_4335(
      {stage015[133], stage015[134], stage015[135], stage015[136], stage015[137]},
      {stage016[153]},
      {stage017[134], stage017[135], stage017[136], stage017[137], stage017[138], stage017[139]},
      {stage019[189], stage018[194], stage017[224], stage016[225], stage015[212]}
   );
   gpc615_5 gpc615_5_4336(
      {stage015[138], stage015[139], stage015[140], stage015[141], stage015[142]},
      {stage016[154]},
      {stage017[140], stage017[141], stage017[142], stage017[143], stage017[144], stage017[145]},
      {stage019[190], stage018[195], stage017[225], stage016[226], stage015[213]}
   );
   gpc615_5 gpc615_5_4337(
      {stage015[143], stage015[144], stage015[145], stage015[146], stage015[147]},
      {stage016[155]},
      {stage017[146], stage017[147], stage017[148], stage017[149], stage017[150], stage017[151]},
      {stage019[191], stage018[196], stage017[226], stage016[227], stage015[214]}
   );
   gpc615_5 gpc615_5_4338(
      {stage015[148], stage015[149], stage015[150], stage015[151], stage015[152]},
      {stage016[156]},
      {stage017[152], stage017[153], stage017[154], stage017[155], stage017[156], stage017[157]},
      {stage019[192], stage018[197], stage017[227], stage016[228], stage015[215]}
   );
   gpc615_5 gpc615_5_4339(
      {stage015[153], stage015[154], stage015[155], stage015[156], stage015[157]},
      {stage016[157]},
      {stage017[158], stage017[159], stage017[160], stage017[161], stage017[162], stage017[163]},
      {stage019[193], stage018[198], stage017[228], stage016[229], stage015[216]}
   );
   gpc615_5 gpc615_5_4340(
      {stage015[158], stage015[159], stage015[160], stage015[161], stage015[162]},
      {stage016[158]},
      {stage017[164], stage017[165], stage017[166], stage017[167], stage017[168], stage017[169]},
      {stage019[194], stage018[199], stage017[229], stage016[230], stage015[217]}
   );
   gpc615_5 gpc615_5_4341(
      {stage015[163], stage015[164], stage015[165], stage015[166], stage015[167]},
      {stage016[159]},
      {stage017[170], stage017[171], stage017[172], stage017[173], stage017[174], stage017[175]},
      {stage019[195], stage018[200], stage017[230], stage016[231], stage015[218]}
   );
   gpc615_5 gpc615_5_4342(
      {stage015[168], stage015[169], stage015[170], stage015[171], stage015[172]},
      {stage016[160]},
      {stage017[176], stage017[177], stage017[178], stage017[179], stage017[180], stage017[181]},
      {stage019[196], stage018[201], stage017[231], stage016[232], stage015[219]}
   );
   gpc615_5 gpc615_5_4343(
      {stage015[173], stage015[174], stage015[175], stage015[176], stage015[177]},
      {stage016[161]},
      {stage017[182], stage017[183], stage017[184], stage017[185], stage017[186], stage017[187]},
      {stage019[197], stage018[202], stage017[232], stage016[233], stage015[220]}
   );
   gpc615_5 gpc615_5_4344(
      {stage015[178], stage015[179], stage015[180], stage015[181], stage015[182]},
      {stage016[162]},
      {stage017[188], stage017[189], stage017[190], stage017[191], stage017[192], stage017[193]},
      {stage019[198], stage018[203], stage017[233], stage016[234], stage015[221]}
   );
   gpc615_5 gpc615_5_4345(
      {stage015[183], stage015[184], stage015[185], stage015[186], stage015[187]},
      {stage016[163]},
      {stage017[194], stage017[195], stage017[196], stage017[197], stage017[198], stage017[199]},
      {stage019[199], stage018[204], stage017[234], stage016[235], stage015[222]}
   );
   gpc1_1 gpc1_1_4346(
      {stage016[164]},
      {stage016[236]}
   );
   gpc1_1 gpc1_1_4347(
      {stage016[165]},
      {stage016[237]}
   );
   gpc1_1 gpc1_1_4348(
      {stage016[166]},
      {stage016[238]}
   );
   gpc606_5 gpc606_5_4349(
      {stage016[167], stage016[168], stage016[169], stage016[170], stage016[171], stage016[172]},
      {stage018[128], stage018[129], stage018[130], stage018[131], stage018[132], stage018[133]},
      {stage020[184], stage019[200], stage018[205], stage017[235], stage016[239]}
   );
   gpc606_5 gpc606_5_4350(
      {stage016[173], stage016[174], stage016[175], stage016[176], stage016[177], stage016[178]},
      {stage018[134], stage018[135], stage018[136], stage018[137], stage018[138], stage018[139]},
      {stage020[185], stage019[201], stage018[206], stage017[236], stage016[240]}
   );
   gpc606_5 gpc606_5_4351(
      {stage016[179], stage016[180], stage016[181], stage016[182], stage016[183], stage016[184]},
      {stage018[140], stage018[141], stage018[142], stage018[143], stage018[144], stage018[145]},
      {stage020[186], stage019[202], stage018[207], stage017[237], stage016[241]}
   );
   gpc606_5 gpc606_5_4352(
      {stage016[185], stage016[186], stage016[187], stage016[188], stage016[189], stage016[190]},
      {stage018[146], stage018[147], stage018[148], stage018[149], stage018[150], stage018[151]},
      {stage020[187], stage019[203], stage018[208], stage017[238], stage016[242]}
   );
   gpc606_5 gpc606_5_4353(
      {stage016[191], stage016[192], stage016[193], stage016[194], stage016[195], stage016[196]},
      {stage018[152], stage018[153], stage018[154], stage018[155], stage018[156], stage018[157]},
      {stage020[188], stage019[204], stage018[209], stage017[239], stage016[243]}
   );
   gpc606_5 gpc606_5_4354(
      {stage016[197], stage016[198], stage016[199], stage016[200], stage016[201], stage016[202]},
      {stage018[158], stage018[159], stage018[160], stage018[161], stage018[162], stage018[163]},
      {stage020[189], stage019[205], stage018[210], stage017[240], stage016[244]}
   );
   gpc1406_5 gpc1406_5_4355(
      {stage016[203], stage016[204], stage016[205], stage016[206], stage016[207], stage016[208]},
      {stage018[164], stage018[165], stage018[166], stage018[167]},
      {stage019[128]},
      {stage020[190], stage019[206], stage018[211], stage017[241], stage016[245]}
   );
   gpc1_1 gpc1_1_4356(
      {stage017[200]},
      {stage017[242]}
   );
   gpc1_1 gpc1_1_4357(
      {stage017[201]},
      {stage017[243]}
   );
   gpc1_1 gpc1_1_4358(
      {stage017[202]},
      {stage017[244]}
   );
   gpc1_1 gpc1_1_4359(
      {stage017[203]},
      {stage017[245]}
   );
   gpc1_1 gpc1_1_4360(
      {stage017[204]},
      {stage017[246]}
   );
   gpc1_1 gpc1_1_4361(
      {stage017[205]},
      {stage017[247]}
   );
   gpc1_1 gpc1_1_4362(
      {stage017[206]},
      {stage017[248]}
   );
   gpc1406_5 gpc1406_5_4363(
      {stage017[207], stage017[208], stage017[209], stage017[210], stage017[211], stage017[212]},
      {stage019[129], stage019[130], stage019[131], stage019[132]},
      {stage020[128]},
      {stage021[201], stage020[191], stage019[207], stage018[212], stage017[249]}
   );
   gpc1406_5 gpc1406_5_4364(
      {stage017[213], stage017[214], stage017[215], stage017[216], stage017[217], stage017[218]},
      {stage019[133], stage019[134], stage019[135], stage019[136]},
      {stage020[129]},
      {stage021[202], stage020[192], stage019[208], stage018[213], stage017[250]}
   );
   gpc1_1 gpc1_1_4365(
      {stage018[168]},
      {stage018[214]}
   );
   gpc1_1 gpc1_1_4366(
      {stage018[169]},
      {stage018[215]}
   );
   gpc1_1 gpc1_1_4367(
      {stage018[170]},
      {stage018[216]}
   );
   gpc1_1 gpc1_1_4368(
      {stage018[171]},
      {stage018[217]}
   );
   gpc1_1 gpc1_1_4369(
      {stage018[172]},
      {stage018[218]}
   );
   gpc615_5 gpc615_5_4370(
      {stage018[173], stage018[174], stage018[175], stage018[176], stage018[177]},
      {stage019[137]},
      {stage020[130], stage020[131], stage020[132], stage020[133], stage020[134], stage020[135]},
      {stage022[180], stage021[203], stage020[193], stage019[209], stage018[219]}
   );
   gpc1406_5 gpc1406_5_4371(
      {stage018[178], stage018[179], stage018[180], stage018[181], stage018[182], stage018[183]},
      {stage020[136], stage020[137], stage020[138], stage020[139]},
      {stage021[128]},
      {stage022[181], stage021[204], stage020[194], stage019[210], stage018[220]}
   );
   gpc135_4 gpc135_4_4372(
      {stage018[184], stage018[185], stage018[186], stage018[187], stage018[188]},
      {stage019[138], stage019[139], stage019[140]},
      {stage020[140]},
      {stage021[205], stage020[195], stage019[211], stage018[221]}
   );
   gpc1_1 gpc1_1_4373(
      {stage019[141]},
      {stage019[212]}
   );
   gpc606_5 gpc606_5_4374(
      {stage019[142], stage019[143], stage019[144], stage019[145], stage019[146], stage019[147]},
      {stage021[129], stage021[130], stage021[131], stage021[132], stage021[133], stage021[134]},
      {stage023[223], stage022[182], stage021[206], stage020[196], stage019[213]}
   );
   gpc615_5 gpc615_5_4375(
      {stage019[148], stage019[149], stage019[150], stage019[151], stage019[152]},
      {stage020[141]},
      {stage021[135], stage021[136], stage021[137], stage021[138], stage021[139], stage021[140]},
      {stage023[224], stage022[183], stage021[207], stage020[197], stage019[214]}
   );
   gpc615_5 gpc615_5_4376(
      {stage019[153], stage019[154], stage019[155], stage019[156], stage019[157]},
      {stage020[142]},
      {stage021[141], stage021[142], stage021[143], stage021[144], stage021[145], stage021[146]},
      {stage023[225], stage022[184], stage021[208], stage020[198], stage019[215]}
   );
   gpc615_5 gpc615_5_4377(
      {stage019[158], stage019[159], stage019[160], stage019[161], stage019[162]},
      {stage020[143]},
      {stage021[147], stage021[148], stage021[149], stage021[150], stage021[151], stage021[152]},
      {stage023[226], stage022[185], stage021[209], stage020[199], stage019[216]}
   );
   gpc615_5 gpc615_5_4378(
      {stage019[163], stage019[164], stage019[165], stage019[166], stage019[167]},
      {stage020[144]},
      {stage021[153], stage021[154], stage021[155], stage021[156], stage021[157], stage021[158]},
      {stage023[227], stage022[186], stage021[210], stage020[200], stage019[217]}
   );
   gpc615_5 gpc615_5_4379(
      {stage019[168], stage019[169], stage019[170], stage019[171], stage019[172]},
      {stage020[145]},
      {stage021[159], stage021[160], stage021[161], stage021[162], stage021[163], stage021[164]},
      {stage023[228], stage022[187], stage021[211], stage020[201], stage019[218]}
   );
   gpc615_5 gpc615_5_4380(
      {stage019[173], stage019[174], stage019[175], stage019[176], stage019[177]},
      {stage020[146]},
      {stage021[165], stage021[166], stage021[167], stage021[168], stage021[169], stage021[170]},
      {stage023[229], stage022[188], stage021[212], stage020[202], stage019[219]}
   );
   gpc615_5 gpc615_5_4381(
      {stage019[178], stage019[179], stage019[180], stage019[181], stage019[182]},
      {stage020[147]},
      {stage021[171], stage021[172], stage021[173], stage021[174], stage021[175], stage021[176]},
      {stage023[230], stage022[189], stage021[213], stage020[203], stage019[220]}
   );
   gpc615_5 gpc615_5_4382(
      {stage019[183], stage019[184], stage019[185], stage019[186], stage019[187]},
      {stage020[148]},
      {stage021[177], stage021[178], stage021[179], stage021[180], stage021[181], stage021[182]},
      {stage023[231], stage022[190], stage021[214], stage020[204], stage019[221]}
   );
   gpc606_5 gpc606_5_4383(
      {stage020[149], stage020[150], stage020[151], stage020[152], stage020[153], stage020[154]},
      {stage022[128], stage022[129], stage022[130], stage022[131], stage022[132], stage022[133]},
      {stage024[188], stage023[232], stage022[191], stage021[215], stage020[205]}
   );
   gpc606_5 gpc606_5_4384(
      {stage020[155], stage020[156], stage020[157], stage020[158], stage020[159], stage020[160]},
      {stage022[134], stage022[135], stage022[136], stage022[137], stage022[138], stage022[139]},
      {stage024[189], stage023[233], stage022[192], stage021[216], stage020[206]}
   );
   gpc606_5 gpc606_5_4385(
      {stage020[161], stage020[162], stage020[163], stage020[164], stage020[165], stage020[166]},
      {stage022[140], stage022[141], stage022[142], stage022[143], stage022[144], stage022[145]},
      {stage024[190], stage023[234], stage022[193], stage021[217], stage020[207]}
   );
   gpc606_5 gpc606_5_4386(
      {stage020[167], stage020[168], stage020[169], stage020[170], stage020[171], stage020[172]},
      {stage022[146], stage022[147], stage022[148], stage022[149], stage022[150], stage022[151]},
      {stage024[191], stage023[235], stage022[194], stage021[218], stage020[208]}
   );
   gpc606_5 gpc606_5_4387(
      {stage020[173], stage020[174], stage020[175], stage020[176], stage020[177], stage020[178]},
      {stage022[152], stage022[153], stage022[154], stage022[155], stage022[156], stage022[157]},
      {stage024[192], stage023[236], stage022[195], stage021[219], stage020[209]}
   );
   gpc606_5 gpc606_5_4388(
      {stage020[179], stage020[180], stage020[181], stage020[182], stage020[183], 1'h0},
      {stage022[158], stage022[159], stage022[160], stage022[161], stage022[162], stage022[163]},
      {stage024[193], stage023[237], stage022[196], stage021[220], stage020[210]}
   );
   gpc1_1 gpc1_1_4389(
      {stage021[183]},
      {stage021[221]}
   );
   gpc1_1 gpc1_1_4390(
      {stage021[184]},
      {stage021[222]}
   );
   gpc1_1 gpc1_1_4391(
      {stage021[185]},
      {stage021[223]}
   );
   gpc1_1 gpc1_1_4392(
      {stage021[186]},
      {stage021[224]}
   );
   gpc1_1 gpc1_1_4393(
      {stage021[187]},
      {stage021[225]}
   );
   gpc1_1 gpc1_1_4394(
      {stage021[188]},
      {stage021[226]}
   );
   gpc1_1 gpc1_1_4395(
      {stage021[189]},
      {stage021[227]}
   );
   gpc1_1 gpc1_1_4396(
      {stage021[190]},
      {stage021[228]}
   );
   gpc1_1 gpc1_1_4397(
      {stage021[191]},
      {stage021[229]}
   );
   gpc1_1 gpc1_1_4398(
      {stage021[192]},
      {stage021[230]}
   );
   gpc1_1 gpc1_1_4399(
      {stage021[193]},
      {stage021[231]}
   );
   gpc1_1 gpc1_1_4400(
      {stage021[194]},
      {stage021[232]}
   );
   gpc1_1 gpc1_1_4401(
      {stage021[195]},
      {stage021[233]}
   );
   gpc1_1 gpc1_1_4402(
      {stage021[196]},
      {stage021[234]}
   );
   gpc1_1 gpc1_1_4403(
      {stage021[197]},
      {stage021[235]}
   );
   gpc1_1 gpc1_1_4404(
      {stage021[198]},
      {stage021[236]}
   );
   gpc1_1 gpc1_1_4405(
      {stage021[199]},
      {stage021[237]}
   );
   gpc1_1 gpc1_1_4406(
      {stage021[200]},
      {stage021[238]}
   );
   gpc1_1 gpc1_1_4407(
      {stage022[164]},
      {stage022[197]}
   );
   gpc1_1 gpc1_1_4408(
      {stage022[165]},
      {stage022[198]}
   );
   gpc7_3 gpc7_3_4409(
      {stage022[166], stage022[167], stage022[168], stage022[169], stage022[170], stage022[171], stage022[172]},
      {stage024[194], stage023[238], stage022[199]}
   );
   gpc7_3 gpc7_3_4410(
      {stage022[173], stage022[174], stage022[175], stage022[176], stage022[177], stage022[178], stage022[179]},
      {stage024[195], stage023[239], stage022[200]}
   );
   gpc1_1 gpc1_1_4411(
      {stage023[128]},
      {stage023[240]}
   );
   gpc1_1 gpc1_1_4412(
      {stage023[129]},
      {stage023[241]}
   );
   gpc1_1 gpc1_1_4413(
      {stage023[130]},
      {stage023[242]}
   );
   gpc1_1 gpc1_1_4414(
      {stage023[131]},
      {stage023[243]}
   );
   gpc1_1 gpc1_1_4415(
      {stage023[132]},
      {stage023[244]}
   );
   gpc1_1 gpc1_1_4416(
      {stage023[133]},
      {stage023[245]}
   );
   gpc1_1 gpc1_1_4417(
      {stage023[134]},
      {stage023[246]}
   );
   gpc1_1 gpc1_1_4418(
      {stage023[135]},
      {stage023[247]}
   );
   gpc1_1 gpc1_1_4419(
      {stage023[136]},
      {stage023[248]}
   );
   gpc1_1 gpc1_1_4420(
      {stage023[137]},
      {stage023[249]}
   );
   gpc1_1 gpc1_1_4421(
      {stage023[138]},
      {stage023[250]}
   );
   gpc606_5 gpc606_5_4422(
      {stage023[139], stage023[140], stage023[141], stage023[142], stage023[143], stage023[144]},
      {stage025[128], stage025[129], stage025[130], stage025[131], stage025[132], stage025[133]},
      {stage027[176], stage026[191], stage025[224], stage024[196], stage023[251]}
   );
   gpc606_5 gpc606_5_4423(
      {stage023[145], stage023[146], stage023[147], stage023[148], stage023[149], stage023[150]},
      {stage025[134], stage025[135], stage025[136], stage025[137], stage025[138], stage025[139]},
      {stage027[177], stage026[192], stage025[225], stage024[197], stage023[252]}
   );
   gpc606_5 gpc606_5_4424(
      {stage023[151], stage023[152], stage023[153], stage023[154], stage023[155], stage023[156]},
      {stage025[140], stage025[141], stage025[142], stage025[143], stage025[144], stage025[145]},
      {stage027[178], stage026[193], stage025[226], stage024[198], stage023[253]}
   );
   gpc606_5 gpc606_5_4425(
      {stage023[157], stage023[158], stage023[159], stage023[160], stage023[161], stage023[162]},
      {stage025[146], stage025[147], stage025[148], stage025[149], stage025[150], stage025[151]},
      {stage027[179], stage026[194], stage025[227], stage024[199], stage023[254]}
   );
   gpc606_5 gpc606_5_4426(
      {stage023[163], stage023[164], stage023[165], stage023[166], stage023[167], stage023[168]},
      {stage025[152], stage025[153], stage025[154], stage025[155], stage025[156], stage025[157]},
      {stage027[180], stage026[195], stage025[228], stage024[200], stage023[255]}
   );
   gpc606_5 gpc606_5_4427(
      {stage023[169], stage023[170], stage023[171], stage023[172], stage023[173], stage023[174]},
      {stage025[158], stage025[159], stage025[160], stage025[161], stage025[162], stage025[163]},
      {stage027[181], stage026[196], stage025[229], stage024[201], stage023[256]}
   );
   gpc606_5 gpc606_5_4428(
      {stage023[175], stage023[176], stage023[177], stage023[178], stage023[179], stage023[180]},
      {stage025[164], stage025[165], stage025[166], stage025[167], stage025[168], stage025[169]},
      {stage027[182], stage026[197], stage025[230], stage024[202], stage023[257]}
   );
   gpc606_5 gpc606_5_4429(
      {stage023[181], stage023[182], stage023[183], stage023[184], stage023[185], stage023[186]},
      {stage025[170], stage025[171], stage025[172], stage025[173], stage025[174], stage025[175]},
      {stage027[183], stage026[198], stage025[231], stage024[203], stage023[258]}
   );
   gpc606_5 gpc606_5_4430(
      {stage023[187], stage023[188], stage023[189], stage023[190], stage023[191], stage023[192]},
      {stage025[176], stage025[177], stage025[178], stage025[179], stage025[180], stage025[181]},
      {stage027[184], stage026[199], stage025[232], stage024[204], stage023[259]}
   );
   gpc606_5 gpc606_5_4431(
      {stage023[193], stage023[194], stage023[195], stage023[196], stage023[197], stage023[198]},
      {stage025[182], stage025[183], stage025[184], stage025[185], stage025[186], stage025[187]},
      {stage027[185], stage026[200], stage025[233], stage024[205], stage023[260]}
   );
   gpc606_5 gpc606_5_4432(
      {stage023[199], stage023[200], stage023[201], stage023[202], stage023[203], stage023[204]},
      {stage025[188], stage025[189], stage025[190], stage025[191], stage025[192], stage025[193]},
      {stage027[186], stage026[201], stage025[234], stage024[206], stage023[261]}
   );
   gpc606_5 gpc606_5_4433(
      {stage023[205], stage023[206], stage023[207], stage023[208], stage023[209], stage023[210]},
      {stage025[194], stage025[195], stage025[196], stage025[197], stage025[198], stage025[199]},
      {stage027[187], stage026[202], stage025[235], stage024[207], stage023[262]}
   );
   gpc606_5 gpc606_5_4434(
      {stage023[211], stage023[212], stage023[213], stage023[214], stage023[215], stage023[216]},
      {stage025[200], stage025[201], stage025[202], stage025[203], stage025[204], stage025[205]},
      {stage027[188], stage026[203], stage025[236], stage024[208], stage023[263]}
   );
   gpc606_5 gpc606_5_4435(
      {stage023[217], stage023[218], stage023[219], stage023[220], stage023[221], stage023[222]},
      {stage025[206], stage025[207], stage025[208], stage025[209], stage025[210], stage025[211]},
      {stage027[189], stage026[204], stage025[237], stage024[209], stage023[264]}
   );
   gpc1_1 gpc1_1_4436(
      {stage024[128]},
      {stage024[210]}
   );
   gpc1_1 gpc1_1_4437(
      {stage024[129]},
      {stage024[211]}
   );
   gpc1_1 gpc1_1_4438(
      {stage024[130]},
      {stage024[212]}
   );
   gpc1_1 gpc1_1_4439(
      {stage024[131]},
      {stage024[213]}
   );
   gpc1_1 gpc1_1_4440(
      {stage024[132]},
      {stage024[214]}
   );
   gpc1_1 gpc1_1_4441(
      {stage024[133]},
      {stage024[215]}
   );
   gpc606_5 gpc606_5_4442(
      {stage024[134], stage024[135], stage024[136], stage024[137], stage024[138], stage024[139]},
      {stage026[128], stage026[129], stage026[130], stage026[131], stage026[132], stage026[133]},
      {stage028[182], stage027[190], stage026[205], stage025[238], stage024[216]}
   );
   gpc606_5 gpc606_5_4443(
      {stage024[140], stage024[141], stage024[142], stage024[143], stage024[144], stage024[145]},
      {stage026[134], stage026[135], stage026[136], stage026[137], stage026[138], stage026[139]},
      {stage028[183], stage027[191], stage026[206], stage025[239], stage024[217]}
   );
   gpc606_5 gpc606_5_4444(
      {stage024[146], stage024[147], stage024[148], stage024[149], stage024[150], stage024[151]},
      {stage026[140], stage026[141], stage026[142], stage026[143], stage026[144], stage026[145]},
      {stage028[184], stage027[192], stage026[207], stage025[240], stage024[218]}
   );
   gpc606_5 gpc606_5_4445(
      {stage024[152], stage024[153], stage024[154], stage024[155], stage024[156], stage024[157]},
      {stage026[146], stage026[147], stage026[148], stage026[149], stage026[150], stage026[151]},
      {stage028[185], stage027[193], stage026[208], stage025[241], stage024[219]}
   );
   gpc606_5 gpc606_5_4446(
      {stage024[158], stage024[159], stage024[160], stage024[161], stage024[162], stage024[163]},
      {stage026[152], stage026[153], stage026[154], stage026[155], stage026[156], stage026[157]},
      {stage028[186], stage027[194], stage026[209], stage025[242], stage024[220]}
   );
   gpc606_5 gpc606_5_4447(
      {stage024[164], stage024[165], stage024[166], stage024[167], stage024[168], stage024[169]},
      {stage026[158], stage026[159], stage026[160], stage026[161], stage026[162], stage026[163]},
      {stage028[187], stage027[195], stage026[210], stage025[243], stage024[221]}
   );
   gpc606_5 gpc606_5_4448(
      {stage024[170], stage024[171], stage024[172], stage024[173], stage024[174], stage024[175]},
      {stage026[164], stage026[165], stage026[166], stage026[167], stage026[168], stage026[169]},
      {stage028[188], stage027[196], stage026[211], stage025[244], stage024[222]}
   );
   gpc606_5 gpc606_5_4449(
      {stage024[176], stage024[177], stage024[178], stage024[179], stage024[180], stage024[181]},
      {stage026[170], stage026[171], stage026[172], stage026[173], stage026[174], stage026[175]},
      {stage028[189], stage027[197], stage026[212], stage025[245], stage024[223]}
   );
   gpc606_5 gpc606_5_4450(
      {stage024[182], stage024[183], stage024[184], stage024[185], stage024[186], stage024[187]},
      {stage026[176], stage026[177], stage026[178], stage026[179], stage026[180], stage026[181]},
      {stage028[190], stage027[198], stage026[213], stage025[246], stage024[224]}
   );
   gpc1_1 gpc1_1_4451(
      {stage025[212]},
      {stage025[247]}
   );
   gpc1_1 gpc1_1_4452(
      {stage025[213]},
      {stage025[248]}
   );
   gpc1_1 gpc1_1_4453(
      {stage025[214]},
      {stage025[249]}
   );
   gpc1_1 gpc1_1_4454(
      {stage025[215]},
      {stage025[250]}
   );
   gpc1_1 gpc1_1_4455(
      {stage025[216]},
      {stage025[251]}
   );
   gpc1_1 gpc1_1_4456(
      {stage025[217]},
      {stage025[252]}
   );
   gpc1_1 gpc1_1_4457(
      {stage025[218]},
      {stage025[253]}
   );
   gpc1_1 gpc1_1_4458(
      {stage025[219]},
      {stage025[254]}
   );
   gpc1_1 gpc1_1_4459(
      {stage025[220]},
      {stage025[255]}
   );
   gpc623_5 gpc623_5_4460(
      {stage025[221], stage025[222], stage025[223]},
      {stage026[182], stage026[183]},
      {stage027[128], stage027[129], stage027[130], stage027[131], stage027[132], stage027[133]},
      {stage029[204], stage028[191], stage027[199], stage026[214], stage025[256]}
   );
   gpc1_1 gpc1_1_4461(
      {stage026[184]},
      {stage026[215]}
   );
   gpc1_1 gpc1_1_4462(
      {stage026[185]},
      {stage026[216]}
   );
   gpc1_1 gpc1_1_4463(
      {stage026[186]},
      {stage026[217]}
   );
   gpc1_1 gpc1_1_4464(
      {stage026[187]},
      {stage026[218]}
   );
   gpc1_1 gpc1_1_4465(
      {stage026[188]},
      {stage026[219]}
   );
   gpc1_1 gpc1_1_4466(
      {stage026[189]},
      {stage026[220]}
   );
   gpc1_1 gpc1_1_4467(
      {stage026[190]},
      {stage026[221]}
   );
   gpc1_1 gpc1_1_4468(
      {stage027[134]},
      {stage027[200]}
   );
   gpc1_1 gpc1_1_4469(
      {stage027[135]},
      {stage027[201]}
   );
   gpc1_1 gpc1_1_4470(
      {stage027[136]},
      {stage027[202]}
   );
   gpc1_1 gpc1_1_4471(
      {stage027[137]},
      {stage027[203]}
   );
   gpc606_5 gpc606_5_4472(
      {stage027[138], stage027[139], stage027[140], stage027[141], stage027[142], stage027[143]},
      {stage029[128], stage029[129], stage029[130], stage029[131], stage029[132], stage029[133]},
      {stage031[171], stage030[184], stage029[205], stage028[192], stage027[204]}
   );
   gpc606_5 gpc606_5_4473(
      {stage027[144], stage027[145], stage027[146], stage027[147], stage027[148], stage027[149]},
      {stage029[134], stage029[135], stage029[136], stage029[137], stage029[138], stage029[139]},
      {stage031[172], stage030[185], stage029[206], stage028[193], stage027[205]}
   );
   gpc606_5 gpc606_5_4474(
      {stage027[150], stage027[151], stage027[152], stage027[153], stage027[154], stage027[155]},
      {stage029[140], stage029[141], stage029[142], stage029[143], stage029[144], stage029[145]},
      {stage031[173], stage030[186], stage029[207], stage028[194], stage027[206]}
   );
   gpc615_5 gpc615_5_4475(
      {stage027[156], stage027[157], stage027[158], stage027[159], stage027[160]},
      {stage028[128]},
      {stage029[146], stage029[147], stage029[148], stage029[149], stage029[150], stage029[151]},
      {stage031[174], stage030[187], stage029[208], stage028[195], stage027[207]}
   );
   gpc615_5 gpc615_5_4476(
      {stage027[161], stage027[162], stage027[163], stage027[164], stage027[165]},
      {stage028[129]},
      {stage029[152], stage029[153], stage029[154], stage029[155], stage029[156], stage029[157]},
      {stage031[175], stage030[188], stage029[209], stage028[196], stage027[208]}
   );
   gpc615_5 gpc615_5_4477(
      {stage027[166], stage027[167], stage027[168], stage027[169], stage027[170]},
      {stage028[130]},
      {stage029[158], stage029[159], stage029[160], stage029[161], stage029[162], stage029[163]},
      {stage031[176], stage030[189], stage029[210], stage028[197], stage027[209]}
   );
   gpc615_5 gpc615_5_4478(
      {stage027[171], stage027[172], stage027[173], stage027[174], stage027[175]},
      {stage028[131]},
      {stage029[164], stage029[165], stage029[166], stage029[167], stage029[168], stage029[169]},
      {stage031[177], stage030[190], stage029[211], stage028[198], stage027[210]}
   );
   gpc1_1 gpc1_1_4479(
      {stage028[132]},
      {stage028[199]}
   );
   gpc1_1 gpc1_1_4480(
      {stage028[133]},
      {stage028[200]}
   );
   gpc1_1 gpc1_1_4481(
      {stage028[134]},
      {stage028[201]}
   );
   gpc1_1 gpc1_1_4482(
      {stage028[135]},
      {stage028[202]}
   );
   gpc1_1 gpc1_1_4483(
      {stage028[136]},
      {stage028[203]}
   );
   gpc1_1 gpc1_1_4484(
      {stage028[137]},
      {stage028[204]}
   );
   gpc1_1 gpc1_1_4485(
      {stage028[138]},
      {stage028[205]}
   );
   gpc1_1 gpc1_1_4486(
      {stage028[139]},
      {stage028[206]}
   );
   gpc1_1 gpc1_1_4487(
      {stage028[140]},
      {stage028[207]}
   );
   gpc1_1 gpc1_1_4488(
      {stage028[141]},
      {stage028[208]}
   );
   gpc1_1 gpc1_1_4489(
      {stage028[142]},
      {stage028[209]}
   );
   gpc1_1 gpc1_1_4490(
      {stage028[143]},
      {stage028[210]}
   );
   gpc1_1 gpc1_1_4491(
      {stage028[144]},
      {stage028[211]}
   );
   gpc1_1 gpc1_1_4492(
      {stage028[145]},
      {stage028[212]}
   );
   gpc1_1 gpc1_1_4493(
      {stage028[146]},
      {stage028[213]}
   );
   gpc1_1 gpc1_1_4494(
      {stage028[147]},
      {stage028[214]}
   );
   gpc1_1 gpc1_1_4495(
      {stage028[148]},
      {stage028[215]}
   );
   gpc1_1 gpc1_1_4496(
      {stage028[149]},
      {stage028[216]}
   );
   gpc1_1 gpc1_1_4497(
      {stage028[150]},
      {stage028[217]}
   );
   gpc1_1 gpc1_1_4498(
      {stage028[151]},
      {stage028[218]}
   );
   gpc606_5 gpc606_5_4499(
      {stage028[152], stage028[153], stage028[154], stage028[155], stage028[156], stage028[157]},
      {stage030[128], stage030[129], stage030[130], stage030[131], stage030[132], stage030[133]},
      {stage032[223], stage031[178], stage030[191], stage029[212], stage028[219]}
   );
   gpc606_5 gpc606_5_4500(
      {stage028[158], stage028[159], stage028[160], stage028[161], stage028[162], stage028[163]},
      {stage030[134], stage030[135], stage030[136], stage030[137], stage030[138], stage030[139]},
      {stage032[224], stage031[179], stage030[192], stage029[213], stage028[220]}
   );
   gpc606_5 gpc606_5_4501(
      {stage028[164], stage028[165], stage028[166], stage028[167], stage028[168], stage028[169]},
      {stage030[140], stage030[141], stage030[142], stage030[143], stage030[144], stage030[145]},
      {stage032[225], stage031[180], stage030[193], stage029[214], stage028[221]}
   );
   gpc606_5 gpc606_5_4502(
      {stage028[170], stage028[171], stage028[172], stage028[173], stage028[174], stage028[175]},
      {stage030[146], stage030[147], stage030[148], stage030[149], stage030[150], stage030[151]},
      {stage032[226], stage031[181], stage030[194], stage029[215], stage028[222]}
   );
   gpc606_5 gpc606_5_4503(
      {stage028[176], stage028[177], stage028[178], stage028[179], stage028[180], stage028[181]},
      {stage030[152], stage030[153], stage030[154], stage030[155], stage030[156], stage030[157]},
      {stage032[227], stage031[182], stage030[195], stage029[216], stage028[223]}
   );
   gpc1_1 gpc1_1_4504(
      {stage029[170]},
      {stage029[217]}
   );
   gpc1_1 gpc1_1_4505(
      {stage029[171]},
      {stage029[218]}
   );
   gpc1_1 gpc1_1_4506(
      {stage029[172]},
      {stage029[219]}
   );
   gpc1_1 gpc1_1_4507(
      {stage029[173]},
      {stage029[220]}
   );
   gpc1_1 gpc1_1_4508(
      {stage029[174]},
      {stage029[221]}
   );
   gpc1_1 gpc1_1_4509(
      {stage029[175]},
      {stage029[222]}
   );
   gpc1_1 gpc1_1_4510(
      {stage029[176]},
      {stage029[223]}
   );
   gpc1_1 gpc1_1_4511(
      {stage029[177]},
      {stage029[224]}
   );
   gpc1_1 gpc1_1_4512(
      {stage029[178]},
      {stage029[225]}
   );
   gpc1_1 gpc1_1_4513(
      {stage029[179]},
      {stage029[226]}
   );
   gpc1_1 gpc1_1_4514(
      {stage029[180]},
      {stage029[227]}
   );
   gpc1_1 gpc1_1_4515(
      {stage029[181]},
      {stage029[228]}
   );
   gpc1_1 gpc1_1_4516(
      {stage029[182]},
      {stage029[229]}
   );
   gpc1_1 gpc1_1_4517(
      {stage029[183]},
      {stage029[230]}
   );
   gpc1_1 gpc1_1_4518(
      {stage029[184]},
      {stage029[231]}
   );
   gpc1_1 gpc1_1_4519(
      {stage029[185]},
      {stage029[232]}
   );
   gpc1_1 gpc1_1_4520(
      {stage029[186]},
      {stage029[233]}
   );
   gpc1_1 gpc1_1_4521(
      {stage029[187]},
      {stage029[234]}
   );
   gpc1_1 gpc1_1_4522(
      {stage029[188]},
      {stage029[235]}
   );
   gpc1_1 gpc1_1_4523(
      {stage029[189]},
      {stage029[236]}
   );
   gpc1_1 gpc1_1_4524(
      {stage029[190]},
      {stage029[237]}
   );
   gpc1_1 gpc1_1_4525(
      {stage029[191]},
      {stage029[238]}
   );
   gpc1_1 gpc1_1_4526(
      {stage029[192]},
      {stage029[239]}
   );
   gpc1_1 gpc1_1_4527(
      {stage029[193]},
      {stage029[240]}
   );
   gpc1_1 gpc1_1_4528(
      {stage029[194]},
      {stage029[241]}
   );
   gpc1_1 gpc1_1_4529(
      {stage029[195]},
      {stage029[242]}
   );
   gpc1_1 gpc1_1_4530(
      {stage029[196]},
      {stage029[243]}
   );
   gpc1_1 gpc1_1_4531(
      {stage029[197]},
      {stage029[244]}
   );
   gpc1_1 gpc1_1_4532(
      {stage029[198]},
      {stage029[245]}
   );
   gpc1_1 gpc1_1_4533(
      {stage029[199]},
      {stage029[246]}
   );
   gpc1_1 gpc1_1_4534(
      {stage029[200]},
      {stage029[247]}
   );
   gpc1_1 gpc1_1_4535(
      {stage029[201]},
      {stage029[248]}
   );
   gpc1_1 gpc1_1_4536(
      {stage029[202]},
      {stage029[249]}
   );
   gpc1_1 gpc1_1_4537(
      {stage029[203]},
      {stage029[250]}
   );
   gpc1_1 gpc1_1_4538(
      {stage030[158]},
      {stage030[196]}
   );
   gpc1_1 gpc1_1_4539(
      {stage030[159]},
      {stage030[197]}
   );
   gpc1_1 gpc1_1_4540(
      {stage030[160]},
      {stage030[198]}
   );
   gpc1_1 gpc1_1_4541(
      {stage030[161]},
      {stage030[199]}
   );
   gpc1_1 gpc1_1_4542(
      {stage030[162]},
      {stage030[200]}
   );
   gpc1_1 gpc1_1_4543(
      {stage030[163]},
      {stage030[201]}
   );
   gpc1_1 gpc1_1_4544(
      {stage030[164]},
      {stage030[202]}
   );
   gpc1_1 gpc1_1_4545(
      {stage030[165]},
      {stage030[203]}
   );
   gpc1_1 gpc1_1_4546(
      {stage030[166]},
      {stage030[204]}
   );
   gpc1_1 gpc1_1_4547(
      {stage030[167]},
      {stage030[205]}
   );
   gpc1_1 gpc1_1_4548(
      {stage030[168]},
      {stage030[206]}
   );
   gpc615_5 gpc615_5_4549(
      {stage030[169], stage030[170], stage030[171], stage030[172], stage030[173]},
      {stage031[128]},
      {stage032[128], stage032[129], stage032[130], stage032[131], stage032[132], stage032[133]},
      {stage034[211], stage033[216], stage032[228], stage031[183], stage030[207]}
   );
   gpc615_5 gpc615_5_4550(
      {stage030[174], stage030[175], stage030[176], stage030[177], stage030[178]},
      {stage031[129]},
      {stage032[134], stage032[135], stage032[136], stage032[137], stage032[138], stage032[139]},
      {stage034[212], stage033[217], stage032[229], stage031[184], stage030[208]}
   );
   gpc615_5 gpc615_5_4551(
      {stage030[179], stage030[180], stage030[181], stage030[182], stage030[183]},
      {stage031[130]},
      {stage032[140], stage032[141], stage032[142], stage032[143], stage032[144], stage032[145]},
      {stage034[213], stage033[218], stage032[230], stage031[185], stage030[209]}
   );
   gpc1_1 gpc1_1_4552(
      {stage031[131]},
      {stage031[186]}
   );
   gpc1_1 gpc1_1_4553(
      {stage031[132]},
      {stage031[187]}
   );
   gpc1_1 gpc1_1_4554(
      {stage031[133]},
      {stage031[188]}
   );
   gpc1_1 gpc1_1_4555(
      {stage031[134]},
      {stage031[189]}
   );
   gpc1_1 gpc1_1_4556(
      {stage031[135]},
      {stage031[190]}
   );
   gpc1_1 gpc1_1_4557(
      {stage031[136]},
      {stage031[191]}
   );
   gpc1_1 gpc1_1_4558(
      {stage031[137]},
      {stage031[192]}
   );
   gpc1_1 gpc1_1_4559(
      {stage031[138]},
      {stage031[193]}
   );
   gpc1_1 gpc1_1_4560(
      {stage031[139]},
      {stage031[194]}
   );
   gpc1_1 gpc1_1_4561(
      {stage031[140]},
      {stage031[195]}
   );
   gpc1_1 gpc1_1_4562(
      {stage031[141]},
      {stage031[196]}
   );
   gpc1_1 gpc1_1_4563(
      {stage031[142]},
      {stage031[197]}
   );
   gpc1_1 gpc1_1_4564(
      {stage031[143]},
      {stage031[198]}
   );
   gpc1_1 gpc1_1_4565(
      {stage031[144]},
      {stage031[199]}
   );
   gpc1_1 gpc1_1_4566(
      {stage031[145]},
      {stage031[200]}
   );
   gpc1_1 gpc1_1_4567(
      {stage031[146]},
      {stage031[201]}
   );
   gpc1_1 gpc1_1_4568(
      {stage031[147]},
      {stage031[202]}
   );
   gpc1_1 gpc1_1_4569(
      {stage031[148]},
      {stage031[203]}
   );
   gpc1_1 gpc1_1_4570(
      {stage031[149]},
      {stage031[204]}
   );
   gpc1_1 gpc1_1_4571(
      {stage031[150]},
      {stage031[205]}
   );
   gpc615_5 gpc615_5_4572(
      {stage031[151], stage031[152], stage031[153], stage031[154], stage031[155]},
      {stage032[146]},
      {stage033[128], stage033[129], stage033[130], stage033[131], stage033[132], stage033[133]},
      {stage035[209], stage034[214], stage033[219], stage032[231], stage031[206]}
   );
   gpc615_5 gpc615_5_4573(
      {stage031[156], stage031[157], stage031[158], stage031[159], stage031[160]},
      {stage032[147]},
      {stage033[134], stage033[135], stage033[136], stage033[137], stage033[138], stage033[139]},
      {stage035[210], stage034[215], stage033[220], stage032[232], stage031[207]}
   );
   gpc615_5 gpc615_5_4574(
      {stage031[161], stage031[162], stage031[163], stage031[164], stage031[165]},
      {stage032[148]},
      {stage033[140], stage033[141], stage033[142], stage033[143], stage033[144], stage033[145]},
      {stage035[211], stage034[216], stage033[221], stage032[233], stage031[208]}
   );
   gpc615_5 gpc615_5_4575(
      {stage031[166], stage031[167], stage031[168], stage031[169], stage031[170]},
      {stage032[149]},
      {stage033[146], stage033[147], stage033[148], stage033[149], stage033[150], stage033[151]},
      {stage035[212], stage034[217], stage033[222], stage032[234], stage031[209]}
   );
   gpc1_1 gpc1_1_4576(
      {stage032[150]},
      {stage032[235]}
   );
   gpc1_1 gpc1_1_4577(
      {stage032[151]},
      {stage032[236]}
   );
   gpc1_1 gpc1_1_4578(
      {stage032[152]},
      {stage032[237]}
   );
   gpc1_1 gpc1_1_4579(
      {stage032[153]},
      {stage032[238]}
   );
   gpc1_1 gpc1_1_4580(
      {stage032[154]},
      {stage032[239]}
   );
   gpc1_1 gpc1_1_4581(
      {stage032[155]},
      {stage032[240]}
   );
   gpc1_1 gpc1_1_4582(
      {stage032[156]},
      {stage032[241]}
   );
   gpc1_1 gpc1_1_4583(
      {stage032[157]},
      {stage032[242]}
   );
   gpc1_1 gpc1_1_4584(
      {stage032[158]},
      {stage032[243]}
   );
   gpc1_1 gpc1_1_4585(
      {stage032[159]},
      {stage032[244]}
   );
   gpc1_1 gpc1_1_4586(
      {stage032[160]},
      {stage032[245]}
   );
   gpc1_1 gpc1_1_4587(
      {stage032[161]},
      {stage032[246]}
   );
   gpc1_1 gpc1_1_4588(
      {stage032[162]},
      {stage032[247]}
   );
   gpc1_1 gpc1_1_4589(
      {stage032[163]},
      {stage032[248]}
   );
   gpc1_1 gpc1_1_4590(
      {stage032[164]},
      {stage032[249]}
   );
   gpc1_1 gpc1_1_4591(
      {stage032[165]},
      {stage032[250]}
   );
   gpc1_1 gpc1_1_4592(
      {stage032[166]},
      {stage032[251]}
   );
   gpc1_1 gpc1_1_4593(
      {stage032[167]},
      {stage032[252]}
   );
   gpc1_1 gpc1_1_4594(
      {stage032[168]},
      {stage032[253]}
   );
   gpc606_5 gpc606_5_4595(
      {stage032[169], stage032[170], stage032[171], stage032[172], stage032[173], stage032[174]},
      {stage034[128], stage034[129], stage034[130], stage034[131], stage034[132], stage034[133]},
      {stage036[173], stage035[213], stage034[218], stage033[223], stage032[254]}
   );
   gpc606_5 gpc606_5_4596(
      {stage032[175], stage032[176], stage032[177], stage032[178], stage032[179], stage032[180]},
      {stage034[134], stage034[135], stage034[136], stage034[137], stage034[138], stage034[139]},
      {stage036[174], stage035[214], stage034[219], stage033[224], stage032[255]}
   );
   gpc606_5 gpc606_5_4597(
      {stage032[181], stage032[182], stage032[183], stage032[184], stage032[185], stage032[186]},
      {stage034[140], stage034[141], stage034[142], stage034[143], stage034[144], stage034[145]},
      {stage036[175], stage035[215], stage034[220], stage033[225], stage032[256]}
   );
   gpc606_5 gpc606_5_4598(
      {stage032[187], stage032[188], stage032[189], stage032[190], stage032[191], stage032[192]},
      {stage034[146], stage034[147], stage034[148], stage034[149], stage034[150], stage034[151]},
      {stage036[176], stage035[216], stage034[221], stage033[226], stage032[257]}
   );
   gpc606_5 gpc606_5_4599(
      {stage032[193], stage032[194], stage032[195], stage032[196], stage032[197], stage032[198]},
      {stage034[152], stage034[153], stage034[154], stage034[155], stage034[156], stage034[157]},
      {stage036[177], stage035[217], stage034[222], stage033[227], stage032[258]}
   );
   gpc606_5 gpc606_5_4600(
      {stage032[199], stage032[200], stage032[201], stage032[202], stage032[203], stage032[204]},
      {stage034[158], stage034[159], stage034[160], stage034[161], stage034[162], stage034[163]},
      {stage036[178], stage035[218], stage034[223], stage033[228], stage032[259]}
   );
   gpc606_5 gpc606_5_4601(
      {stage032[205], stage032[206], stage032[207], stage032[208], stage032[209], stage032[210]},
      {stage034[164], stage034[165], stage034[166], stage034[167], stage034[168], stage034[169]},
      {stage036[179], stage035[219], stage034[224], stage033[229], stage032[260]}
   );
   gpc606_5 gpc606_5_4602(
      {stage032[211], stage032[212], stage032[213], stage032[214], stage032[215], stage032[216]},
      {stage034[170], stage034[171], stage034[172], stage034[173], stage034[174], stage034[175]},
      {stage036[180], stage035[220], stage034[225], stage033[230], stage032[261]}
   );
   gpc606_5 gpc606_5_4603(
      {stage032[217], stage032[218], stage032[219], stage032[220], stage032[221], stage032[222]},
      {stage034[176], stage034[177], stage034[178], stage034[179], stage034[180], stage034[181]},
      {stage036[181], stage035[221], stage034[226], stage033[231], stage032[262]}
   );
   gpc1_1 gpc1_1_4604(
      {stage033[152]},
      {stage033[232]}
   );
   gpc1_1 gpc1_1_4605(
      {stage033[153]},
      {stage033[233]}
   );
   gpc1_1 gpc1_1_4606(
      {stage033[154]},
      {stage033[234]}
   );
   gpc1_1 gpc1_1_4607(
      {stage033[155]},
      {stage033[235]}
   );
   gpc1_1 gpc1_1_4608(
      {stage033[156]},
      {stage033[236]}
   );
   gpc1_1 gpc1_1_4609(
      {stage033[157]},
      {stage033[237]}
   );
   gpc1_1 gpc1_1_4610(
      {stage033[158]},
      {stage033[238]}
   );
   gpc1_1 gpc1_1_4611(
      {stage033[159]},
      {stage033[239]}
   );
   gpc1_1 gpc1_1_4612(
      {stage033[160]},
      {stage033[240]}
   );
   gpc1_1 gpc1_1_4613(
      {stage033[161]},
      {stage033[241]}
   );
   gpc1_1 gpc1_1_4614(
      {stage033[162]},
      {stage033[242]}
   );
   gpc1_1 gpc1_1_4615(
      {stage033[163]},
      {stage033[243]}
   );
   gpc1_1 gpc1_1_4616(
      {stage033[164]},
      {stage033[244]}
   );
   gpc1_1 gpc1_1_4617(
      {stage033[165]},
      {stage033[245]}
   );
   gpc1_1 gpc1_1_4618(
      {stage033[166]},
      {stage033[246]}
   );
   gpc1_1 gpc1_1_4619(
      {stage033[167]},
      {stage033[247]}
   );
   gpc1_1 gpc1_1_4620(
      {stage033[168]},
      {stage033[248]}
   );
   gpc1_1 gpc1_1_4621(
      {stage033[169]},
      {stage033[249]}
   );
   gpc1_1 gpc1_1_4622(
      {stage033[170]},
      {stage033[250]}
   );
   gpc1_1 gpc1_1_4623(
      {stage033[171]},
      {stage033[251]}
   );
   gpc1_1 gpc1_1_4624(
      {stage033[172]},
      {stage033[252]}
   );
   gpc1_1 gpc1_1_4625(
      {stage033[173]},
      {stage033[253]}
   );
   gpc1_1 gpc1_1_4626(
      {stage033[174]},
      {stage033[254]}
   );
   gpc1_1 gpc1_1_4627(
      {stage033[175]},
      {stage033[255]}
   );
   gpc1_1 gpc1_1_4628(
      {stage033[176]},
      {stage033[256]}
   );
   gpc1_1 gpc1_1_4629(
      {stage033[177]},
      {stage033[257]}
   );
   gpc1_1 gpc1_1_4630(
      {stage033[178]},
      {stage033[258]}
   );
   gpc1_1 gpc1_1_4631(
      {stage033[179]},
      {stage033[259]}
   );
   gpc606_5 gpc606_5_4632(
      {stage033[180], stage033[181], stage033[182], stage033[183], stage033[184], stage033[185]},
      {stage035[128], stage035[129], stage035[130], stage035[131], stage035[132], stage035[133]},
      {stage037[200], stage036[182], stage035[222], stage034[227], stage033[260]}
   );
   gpc606_5 gpc606_5_4633(
      {stage033[186], stage033[187], stage033[188], stage033[189], stage033[190], stage033[191]},
      {stage035[134], stage035[135], stage035[136], stage035[137], stage035[138], stage035[139]},
      {stage037[201], stage036[183], stage035[223], stage034[228], stage033[261]}
   );
   gpc606_5 gpc606_5_4634(
      {stage033[192], stage033[193], stage033[194], stage033[195], stage033[196], stage033[197]},
      {stage035[140], stage035[141], stage035[142], stage035[143], stage035[144], stage035[145]},
      {stage037[202], stage036[184], stage035[224], stage034[229], stage033[262]}
   );
   gpc606_5 gpc606_5_4635(
      {stage033[198], stage033[199], stage033[200], stage033[201], stage033[202], stage033[203]},
      {stage035[146], stage035[147], stage035[148], stage035[149], stage035[150], stage035[151]},
      {stage037[203], stage036[185], stage035[225], stage034[230], stage033[263]}
   );
   gpc606_5 gpc606_5_4636(
      {stage033[204], stage033[205], stage033[206], stage033[207], stage033[208], stage033[209]},
      {stage035[152], stage035[153], stage035[154], stage035[155], stage035[156], stage035[157]},
      {stage037[204], stage036[186], stage035[226], stage034[231], stage033[264]}
   );
   gpc606_5 gpc606_5_4637(
      {stage033[210], stage033[211], stage033[212], stage033[213], stage033[214], stage033[215]},
      {stage035[158], stage035[159], stage035[160], stage035[161], stage035[162], stage035[163]},
      {stage037[205], stage036[187], stage035[227], stage034[232], stage033[265]}
   );
   gpc1_1 gpc1_1_4638(
      {stage034[182]},
      {stage034[233]}
   );
   gpc1_1 gpc1_1_4639(
      {stage034[183]},
      {stage034[234]}
   );
   gpc1_1 gpc1_1_4640(
      {stage034[184]},
      {stage034[235]}
   );
   gpc1_1 gpc1_1_4641(
      {stage034[185]},
      {stage034[236]}
   );
   gpc1_1 gpc1_1_4642(
      {stage034[186]},
      {stage034[237]}
   );
   gpc1_1 gpc1_1_4643(
      {stage034[187]},
      {stage034[238]}
   );
   gpc1_1 gpc1_1_4644(
      {stage034[188]},
      {stage034[239]}
   );
   gpc1_1 gpc1_1_4645(
      {stage034[189]},
      {stage034[240]}
   );
   gpc1_1 gpc1_1_4646(
      {stage034[190]},
      {stage034[241]}
   );
   gpc1_1 gpc1_1_4647(
      {stage034[191]},
      {stage034[242]}
   );
   gpc1_1 gpc1_1_4648(
      {stage034[192]},
      {stage034[243]}
   );
   gpc1_1 gpc1_1_4649(
      {stage034[193]},
      {stage034[244]}
   );
   gpc1_1 gpc1_1_4650(
      {stage034[194]},
      {stage034[245]}
   );
   gpc1_1 gpc1_1_4651(
      {stage034[195]},
      {stage034[246]}
   );
   gpc1_1 gpc1_1_4652(
      {stage034[196]},
      {stage034[247]}
   );
   gpc1_1 gpc1_1_4653(
      {stage034[197]},
      {stage034[248]}
   );
   gpc1_1 gpc1_1_4654(
      {stage034[198]},
      {stage034[249]}
   );
   gpc1_1 gpc1_1_4655(
      {stage034[199]},
      {stage034[250]}
   );
   gpc1_1 gpc1_1_4656(
      {stage034[200]},
      {stage034[251]}
   );
   gpc1_1 gpc1_1_4657(
      {stage034[201]},
      {stage034[252]}
   );
   gpc1_1 gpc1_1_4658(
      {stage034[202]},
      {stage034[253]}
   );
   gpc1_1 gpc1_1_4659(
      {stage034[203]},
      {stage034[254]}
   );
   gpc1_1 gpc1_1_4660(
      {stage034[204]},
      {stage034[255]}
   );
   gpc1_1 gpc1_1_4661(
      {stage034[205]},
      {stage034[256]}
   );
   gpc1_1 gpc1_1_4662(
      {stage034[206]},
      {stage034[257]}
   );
   gpc1_1 gpc1_1_4663(
      {stage034[207]},
      {stage034[258]}
   );
   gpc1_1 gpc1_1_4664(
      {stage034[208]},
      {stage034[259]}
   );
   gpc1_1 gpc1_1_4665(
      {stage034[209]},
      {stage034[260]}
   );
   gpc1_1 gpc1_1_4666(
      {stage034[210]},
      {stage034[261]}
   );
   gpc615_5 gpc615_5_4667(
      {stage035[164], stage035[165], stage035[166], stage035[167], stage035[168]},
      {stage036[128]},
      {stage037[128], stage037[129], stage037[130], stage037[131], stage037[132], stage037[133]},
      {stage039[189], stage038[193], stage037[206], stage036[188], stage035[228]}
   );
   gpc615_5 gpc615_5_4668(
      {stage035[169], stage035[170], stage035[171], stage035[172], stage035[173]},
      {stage036[129]},
      {stage037[134], stage037[135], stage037[136], stage037[137], stage037[138], stage037[139]},
      {stage039[190], stage038[194], stage037[207], stage036[189], stage035[229]}
   );
   gpc615_5 gpc615_5_4669(
      {stage035[174], stage035[175], stage035[176], stage035[177], stage035[178]},
      {stage036[130]},
      {stage037[140], stage037[141], stage037[142], stage037[143], stage037[144], stage037[145]},
      {stage039[191], stage038[195], stage037[208], stage036[190], stage035[230]}
   );
   gpc615_5 gpc615_5_4670(
      {stage035[179], stage035[180], stage035[181], stage035[182], stage035[183]},
      {stage036[131]},
      {stage037[146], stage037[147], stage037[148], stage037[149], stage037[150], stage037[151]},
      {stage039[192], stage038[196], stage037[209], stage036[191], stage035[231]}
   );
   gpc615_5 gpc615_5_4671(
      {stage035[184], stage035[185], stage035[186], stage035[187], stage035[188]},
      {stage036[132]},
      {stage037[152], stage037[153], stage037[154], stage037[155], stage037[156], stage037[157]},
      {stage039[193], stage038[197], stage037[210], stage036[192], stage035[232]}
   );
   gpc615_5 gpc615_5_4672(
      {stage035[189], stage035[190], stage035[191], stage035[192], stage035[193]},
      {stage036[133]},
      {stage037[158], stage037[159], stage037[160], stage037[161], stage037[162], stage037[163]},
      {stage039[194], stage038[198], stage037[211], stage036[193], stage035[233]}
   );
   gpc615_5 gpc615_5_4673(
      {stage035[194], stage035[195], stage035[196], stage035[197], stage035[198]},
      {stage036[134]},
      {stage037[164], stage037[165], stage037[166], stage037[167], stage037[168], stage037[169]},
      {stage039[195], stage038[199], stage037[212], stage036[194], stage035[234]}
   );
   gpc615_5 gpc615_5_4674(
      {stage035[199], stage035[200], stage035[201], stage035[202], stage035[203]},
      {stage036[135]},
      {stage037[170], stage037[171], stage037[172], stage037[173], stage037[174], stage037[175]},
      {stage039[196], stage038[200], stage037[213], stage036[195], stage035[235]}
   );
   gpc615_5 gpc615_5_4675(
      {stage035[204], stage035[205], stage035[206], stage035[207], stage035[208]},
      {stage036[136]},
      {stage037[176], stage037[177], stage037[178], stage037[179], stage037[180], stage037[181]},
      {stage039[197], stage038[201], stage037[214], stage036[196], stage035[236]}
   );
   gpc606_5 gpc606_5_4676(
      {stage036[137], stage036[138], stage036[139], stage036[140], stage036[141], stage036[142]},
      {stage038[128], stage038[129], stage038[130], stage038[131], stage038[132], stage038[133]},
      {stage040[218], stage039[198], stage038[202], stage037[215], stage036[197]}
   );
   gpc606_5 gpc606_5_4677(
      {stage036[143], stage036[144], stage036[145], stage036[146], stage036[147], stage036[148]},
      {stage038[134], stage038[135], stage038[136], stage038[137], stage038[138], stage038[139]},
      {stage040[219], stage039[199], stage038[203], stage037[216], stage036[198]}
   );
   gpc606_5 gpc606_5_4678(
      {stage036[149], stage036[150], stage036[151], stage036[152], stage036[153], stage036[154]},
      {stage038[140], stage038[141], stage038[142], stage038[143], stage038[144], stage038[145]},
      {stage040[220], stage039[200], stage038[204], stage037[217], stage036[199]}
   );
   gpc606_5 gpc606_5_4679(
      {stage036[155], stage036[156], stage036[157], stage036[158], stage036[159], stage036[160]},
      {stage038[146], stage038[147], stage038[148], stage038[149], stage038[150], stage038[151]},
      {stage040[221], stage039[201], stage038[205], stage037[218], stage036[200]}
   );
   gpc606_5 gpc606_5_4680(
      {stage036[161], stage036[162], stage036[163], stage036[164], stage036[165], stage036[166]},
      {stage038[152], stage038[153], stage038[154], stage038[155], stage038[156], stage038[157]},
      {stage040[222], stage039[202], stage038[206], stage037[219], stage036[201]}
   );
   gpc606_5 gpc606_5_4681(
      {stage036[167], stage036[168], stage036[169], stage036[170], stage036[171], stage036[172]},
      {stage038[158], stage038[159], stage038[160], stage038[161], stage038[162], stage038[163]},
      {stage040[223], stage039[203], stage038[207], stage037[220], stage036[202]}
   );
   gpc1_1 gpc1_1_4682(
      {stage037[182]},
      {stage037[221]}
   );
   gpc1_1 gpc1_1_4683(
      {stage037[183]},
      {stage037[222]}
   );
   gpc1_1 gpc1_1_4684(
      {stage037[184]},
      {stage037[223]}
   );
   gpc1_1 gpc1_1_4685(
      {stage037[185]},
      {stage037[224]}
   );
   gpc1_1 gpc1_1_4686(
      {stage037[186]},
      {stage037[225]}
   );
   gpc1_1 gpc1_1_4687(
      {stage037[187]},
      {stage037[226]}
   );
   gpc606_5 gpc606_5_4688(
      {stage037[188], stage037[189], stage037[190], stage037[191], stage037[192], stage037[193]},
      {stage039[128], stage039[129], stage039[130], stage039[131], stage039[132], stage039[133]},
      {stage041[202], stage040[224], stage039[204], stage038[208], stage037[227]}
   );
   gpc606_5 gpc606_5_4689(
      {stage037[194], stage037[195], stage037[196], stage037[197], stage037[198], stage037[199]},
      {stage039[134], stage039[135], stage039[136], stage039[137], stage039[138], stage039[139]},
      {stage041[203], stage040[225], stage039[205], stage038[209], stage037[228]}
   );
   gpc1_1 gpc1_1_4690(
      {stage038[164]},
      {stage038[210]}
   );
   gpc1_1 gpc1_1_4691(
      {stage038[165]},
      {stage038[211]}
   );
   gpc1_1 gpc1_1_4692(
      {stage038[166]},
      {stage038[212]}
   );
   gpc1_1 gpc1_1_4693(
      {stage038[167]},
      {stage038[213]}
   );
   gpc1_1 gpc1_1_4694(
      {stage038[168]},
      {stage038[214]}
   );
   gpc1_1 gpc1_1_4695(
      {stage038[169]},
      {stage038[215]}
   );
   gpc1_1 gpc1_1_4696(
      {stage038[170]},
      {stage038[216]}
   );
   gpc1_1 gpc1_1_4697(
      {stage038[171]},
      {stage038[217]}
   );
   gpc1_1 gpc1_1_4698(
      {stage038[172]},
      {stage038[218]}
   );
   gpc615_5 gpc615_5_4699(
      {stage038[173], stage038[174], stage038[175], stage038[176], stage038[177]},
      {stage039[140]},
      {stage040[128], stage040[129], stage040[130], stage040[131], stage040[132], stage040[133]},
      {stage042[209], stage041[204], stage040[226], stage039[206], stage038[219]}
   );
   gpc615_5 gpc615_5_4700(
      {stage038[178], stage038[179], stage038[180], stage038[181], stage038[182]},
      {stage039[141]},
      {stage040[134], stage040[135], stage040[136], stage040[137], stage040[138], stage040[139]},
      {stage042[210], stage041[205], stage040[227], stage039[207], stage038[220]}
   );
   gpc615_5 gpc615_5_4701(
      {stage038[183], stage038[184], stage038[185], stage038[186], stage038[187]},
      {stage039[142]},
      {stage040[140], stage040[141], stage040[142], stage040[143], stage040[144], stage040[145]},
      {stage042[211], stage041[206], stage040[228], stage039[208], stage038[221]}
   );
   gpc615_5 gpc615_5_4702(
      {stage038[188], stage038[189], stage038[190], stage038[191], stage038[192]},
      {stage039[143]},
      {stage040[146], stage040[147], stage040[148], stage040[149], stage040[150], stage040[151]},
      {stage042[212], stage041[207], stage040[229], stage039[209], stage038[222]}
   );
   gpc1_1 gpc1_1_4703(
      {stage039[144]},
      {stage039[210]}
   );
   gpc1_1 gpc1_1_4704(
      {stage039[145]},
      {stage039[211]}
   );
   gpc1_1 gpc1_1_4705(
      {stage039[146]},
      {stage039[212]}
   );
   gpc1_1 gpc1_1_4706(
      {stage039[147]},
      {stage039[213]}
   );
   gpc1_1 gpc1_1_4707(
      {stage039[148]},
      {stage039[214]}
   );
   gpc1_1 gpc1_1_4708(
      {stage039[149]},
      {stage039[215]}
   );
   gpc1_1 gpc1_1_4709(
      {stage039[150]},
      {stage039[216]}
   );
   gpc606_5 gpc606_5_4710(
      {stage039[151], stage039[152], stage039[153], stage039[154], stage039[155], stage039[156]},
      {stage041[128], stage041[129], stage041[130], stage041[131], stage041[132], stage041[133]},
      {stage043[166], stage042[213], stage041[208], stage040[230], stage039[217]}
   );
   gpc606_5 gpc606_5_4711(
      {stage039[157], stage039[158], stage039[159], stage039[160], stage039[161], stage039[162]},
      {stage041[134], stage041[135], stage041[136], stage041[137], stage041[138], stage041[139]},
      {stage043[167], stage042[214], stage041[209], stage040[231], stage039[218]}
   );
   gpc606_5 gpc606_5_4712(
      {stage039[163], stage039[164], stage039[165], stage039[166], stage039[167], stage039[168]},
      {stage041[140], stage041[141], stage041[142], stage041[143], stage041[144], stage041[145]},
      {stage043[168], stage042[215], stage041[210], stage040[232], stage039[219]}
   );
   gpc615_5 gpc615_5_4713(
      {stage039[169], stage039[170], stage039[171], stage039[172], stage039[173]},
      {stage040[152]},
      {stage041[146], stage041[147], stage041[148], stage041[149], stage041[150], stage041[151]},
      {stage043[169], stage042[216], stage041[211], stage040[233], stage039[220]}
   );
   gpc615_5 gpc615_5_4714(
      {stage039[174], stage039[175], stage039[176], stage039[177], stage039[178]},
      {stage040[153]},
      {stage041[152], stage041[153], stage041[154], stage041[155], stage041[156], stage041[157]},
      {stage043[170], stage042[217], stage041[212], stage040[234], stage039[221]}
   );
   gpc615_5 gpc615_5_4715(
      {stage039[179], stage039[180], stage039[181], stage039[182], stage039[183]},
      {stage040[154]},
      {stage041[158], stage041[159], stage041[160], stage041[161], stage041[162], stage041[163]},
      {stage043[171], stage042[218], stage041[213], stage040[235], stage039[222]}
   );
   gpc615_5 gpc615_5_4716(
      {stage039[184], stage039[185], stage039[186], stage039[187], stage039[188]},
      {stage040[155]},
      {stage041[164], stage041[165], stage041[166], stage041[167], stage041[168], stage041[169]},
      {stage043[172], stage042[219], stage041[214], stage040[236], stage039[223]}
   );
   gpc1_1 gpc1_1_4717(
      {stage040[156]},
      {stage040[237]}
   );
   gpc1_1 gpc1_1_4718(
      {stage040[157]},
      {stage040[238]}
   );
   gpc1_1 gpc1_1_4719(
      {stage040[158]},
      {stage040[239]}
   );
   gpc1_1 gpc1_1_4720(
      {stage040[159]},
      {stage040[240]}
   );
   gpc1_1 gpc1_1_4721(
      {stage040[160]},
      {stage040[241]}
   );
   gpc1_1 gpc1_1_4722(
      {stage040[161]},
      {stage040[242]}
   );
   gpc1_1 gpc1_1_4723(
      {stage040[162]},
      {stage040[243]}
   );
   gpc1_1 gpc1_1_4724(
      {stage040[163]},
      {stage040[244]}
   );
   gpc1_1 gpc1_1_4725(
      {stage040[164]},
      {stage040[245]}
   );
   gpc1_1 gpc1_1_4726(
      {stage040[165]},
      {stage040[246]}
   );
   gpc1_1 gpc1_1_4727(
      {stage040[166]},
      {stage040[247]}
   );
   gpc1_1 gpc1_1_4728(
      {stage040[167]},
      {stage040[248]}
   );
   gpc1_1 gpc1_1_4729(
      {stage040[168]},
      {stage040[249]}
   );
   gpc1_1 gpc1_1_4730(
      {stage040[169]},
      {stage040[250]}
   );
   gpc1_1 gpc1_1_4731(
      {stage040[170]},
      {stage040[251]}
   );
   gpc1_1 gpc1_1_4732(
      {stage040[171]},
      {stage040[252]}
   );
   gpc1_1 gpc1_1_4733(
      {stage040[172]},
      {stage040[253]}
   );
   gpc1_1 gpc1_1_4734(
      {stage040[173]},
      {stage040[254]}
   );
   gpc1_1 gpc1_1_4735(
      {stage040[174]},
      {stage040[255]}
   );
   gpc1_1 gpc1_1_4736(
      {stage040[175]},
      {stage040[256]}
   );
   gpc623_5 gpc623_5_4737(
      {stage040[176], stage040[177], stage040[178]},
      {stage041[170], stage041[171]},
      {stage042[128], stage042[129], stage042[130], stage042[131], stage042[132], stage042[133]},
      {stage044[179], stage043[173], stage042[220], stage041[215], stage040[257]}
   );
   gpc623_5 gpc623_5_4738(
      {stage040[179], stage040[180], stage040[181]},
      {stage041[172], stage041[173]},
      {stage042[134], stage042[135], stage042[136], stage042[137], stage042[138], stage042[139]},
      {stage044[180], stage043[174], stage042[221], stage041[216], stage040[258]}
   );
   gpc623_5 gpc623_5_4739(
      {stage040[182], stage040[183], stage040[184]},
      {stage041[174], stage041[175]},
      {stage042[140], stage042[141], stage042[142], stage042[143], stage042[144], stage042[145]},
      {stage044[181], stage043[175], stage042[222], stage041[217], stage040[259]}
   );
   gpc623_5 gpc623_5_4740(
      {stage040[185], stage040[186], stage040[187]},
      {stage041[176], stage041[177]},
      {stage042[146], stage042[147], stage042[148], stage042[149], stage042[150], stage042[151]},
      {stage044[182], stage043[176], stage042[223], stage041[218], stage040[260]}
   );
   gpc623_5 gpc623_5_4741(
      {stage040[188], stage040[189], stage040[190]},
      {stage041[178], stage041[179]},
      {stage042[152], stage042[153], stage042[154], stage042[155], stage042[156], stage042[157]},
      {stage044[183], stage043[177], stage042[224], stage041[219], stage040[261]}
   );
   gpc623_5 gpc623_5_4742(
      {stage040[191], stage040[192], stage040[193]},
      {stage041[180], stage041[181]},
      {stage042[158], stage042[159], stage042[160], stage042[161], stage042[162], stage042[163]},
      {stage044[184], stage043[178], stage042[225], stage041[220], stage040[262]}
   );
   gpc623_5 gpc623_5_4743(
      {stage040[194], stage040[195], stage040[196]},
      {stage041[182], stage041[183]},
      {stage042[164], stage042[165], stage042[166], stage042[167], stage042[168], stage042[169]},
      {stage044[185], stage043[179], stage042[226], stage041[221], stage040[263]}
   );
   gpc623_5 gpc623_5_4744(
      {stage040[197], stage040[198], stage040[199]},
      {stage041[184], stage041[185]},
      {stage042[170], stage042[171], stage042[172], stage042[173], stage042[174], stage042[175]},
      {stage044[186], stage043[180], stage042[227], stage041[222], stage040[264]}
   );
   gpc606_5 gpc606_5_4745(
      {stage040[200], stage040[201], stage040[202], stage040[203], stage040[204], stage040[205]},
      {stage042[176], stage042[177], stage042[178], stage042[179], stage042[180], stage042[181]},
      {stage044[187], stage043[181], stage042[228], stage041[223], stage040[265]}
   );
   gpc606_5 gpc606_5_4746(
      {stage040[206], stage040[207], stage040[208], stage040[209], stage040[210], stage040[211]},
      {stage042[182], stage042[183], stage042[184], stage042[185], stage042[186], stage042[187]},
      {stage044[188], stage043[182], stage042[229], stage041[224], stage040[266]}
   );
   gpc606_5 gpc606_5_4747(
      {stage040[212], stage040[213], stage040[214], stage040[215], stage040[216], stage040[217]},
      {stage042[188], stage042[189], stage042[190], stage042[191], stage042[192], stage042[193]},
      {stage044[189], stage043[183], stage042[230], stage041[225], stage040[267]}
   );
   gpc1_1 gpc1_1_4748(
      {stage041[186]},
      {stage041[226]}
   );
   gpc1_1 gpc1_1_4749(
      {stage041[187]},
      {stage041[227]}
   );
   gpc1_1 gpc1_1_4750(
      {stage041[188]},
      {stage041[228]}
   );
   gpc1_1 gpc1_1_4751(
      {stage041[189]},
      {stage041[229]}
   );
   gpc1_1 gpc1_1_4752(
      {stage041[190]},
      {stage041[230]}
   );
   gpc1_1 gpc1_1_4753(
      {stage041[191]},
      {stage041[231]}
   );
   gpc1_1 gpc1_1_4754(
      {stage041[192]},
      {stage041[232]}
   );
   gpc1_1 gpc1_1_4755(
      {stage041[193]},
      {stage041[233]}
   );
   gpc1_1 gpc1_1_4756(
      {stage041[194]},
      {stage041[234]}
   );
   gpc1_1 gpc1_1_4757(
      {stage041[195]},
      {stage041[235]}
   );
   gpc606_5 gpc606_5_4758(
      {stage041[196], stage041[197], stage041[198], stage041[199], stage041[200], stage041[201]},
      {stage043[128], stage043[129], stage043[130], stage043[131], stage043[132], stage043[133]},
      {stage045[204], stage044[190], stage043[184], stage042[231], stage041[236]}
   );
   gpc1_1 gpc1_1_4759(
      {stage042[194]},
      {stage042[232]}
   );
   gpc1_1 gpc1_1_4760(
      {stage042[195]},
      {stage042[233]}
   );
   gpc1_1 gpc1_1_4761(
      {stage042[196]},
      {stage042[234]}
   );
   gpc1_1 gpc1_1_4762(
      {stage042[197]},
      {stage042[235]}
   );
   gpc1_1 gpc1_1_4763(
      {stage042[198]},
      {stage042[236]}
   );
   gpc1_1 gpc1_1_4764(
      {stage042[199]},
      {stage042[237]}
   );
   gpc1_1 gpc1_1_4765(
      {stage042[200]},
      {stage042[238]}
   );
   gpc1_1 gpc1_1_4766(
      {stage042[201]},
      {stage042[239]}
   );
   gpc1_1 gpc1_1_4767(
      {stage042[202]},
      {stage042[240]}
   );
   gpc1_1 gpc1_1_4768(
      {stage042[203]},
      {stage042[241]}
   );
   gpc1_1 gpc1_1_4769(
      {stage042[204]},
      {stage042[242]}
   );
   gpc1_1 gpc1_1_4770(
      {stage042[205]},
      {stage042[243]}
   );
   gpc1_1 gpc1_1_4771(
      {stage042[206]},
      {stage042[244]}
   );
   gpc1_1 gpc1_1_4772(
      {stage042[207]},
      {stage042[245]}
   );
   gpc1_1 gpc1_1_4773(
      {stage042[208]},
      {stage042[246]}
   );
   gpc1_1 gpc1_1_4774(
      {stage043[134]},
      {stage043[185]}
   );
   gpc1_1 gpc1_1_4775(
      {stage043[135]},
      {stage043[186]}
   );
   gpc1_1 gpc1_1_4776(
      {stage043[136]},
      {stage043[187]}
   );
   gpc1_1 gpc1_1_4777(
      {stage043[137]},
      {stage043[188]}
   );
   gpc1_1 gpc1_1_4778(
      {stage043[138]},
      {stage043[189]}
   );
   gpc1_1 gpc1_1_4779(
      {stage043[139]},
      {stage043[190]}
   );
   gpc606_5 gpc606_5_4780(
      {stage043[140], stage043[141], stage043[142], stage043[143], stage043[144], stage043[145]},
      {stage045[128], stage045[129], stage045[130], stage045[131], stage045[132], stage045[133]},
      {stage047[170], stage046[216], stage045[205], stage044[191], stage043[191]}
   );
   gpc615_5 gpc615_5_4781(
      {stage043[146], stage043[147], stage043[148], stage043[149], stage043[150]},
      {stage044[128]},
      {stage045[134], stage045[135], stage045[136], stage045[137], stage045[138], stage045[139]},
      {stage047[171], stage046[217], stage045[206], stage044[192], stage043[192]}
   );
   gpc615_5 gpc615_5_4782(
      {stage043[151], stage043[152], stage043[153], stage043[154], stage043[155]},
      {stage044[129]},
      {stage045[140], stage045[141], stage045[142], stage045[143], stage045[144], stage045[145]},
      {stage047[172], stage046[218], stage045[207], stage044[193], stage043[193]}
   );
   gpc615_5 gpc615_5_4783(
      {stage043[156], stage043[157], stage043[158], stage043[159], stage043[160]},
      {stage044[130]},
      {stage045[146], stage045[147], stage045[148], stage045[149], stage045[150], stage045[151]},
      {stage047[173], stage046[219], stage045[208], stage044[194], stage043[194]}
   );
   gpc615_5 gpc615_5_4784(
      {stage043[161], stage043[162], stage043[163], stage043[164], stage043[165]},
      {stage044[131]},
      {stage045[152], stage045[153], stage045[154], stage045[155], stage045[156], stage045[157]},
      {stage047[174], stage046[220], stage045[209], stage044[195], stage043[195]}
   );
   gpc623_5 gpc623_5_4785(
      {stage044[132], stage044[133], stage044[134]},
      {stage045[158], stage045[159]},
      {stage046[128], stage046[129], stage046[130], stage046[131], stage046[132], stage046[133]},
      {stage048[230], stage047[175], stage046[221], stage045[210], stage044[196]}
   );
   gpc623_5 gpc623_5_4786(
      {stage044[135], stage044[136], stage044[137]},
      {stage045[160], stage045[161]},
      {stage046[134], stage046[135], stage046[136], stage046[137], stage046[138], stage046[139]},
      {stage048[231], stage047[176], stage046[222], stage045[211], stage044[197]}
   );
   gpc623_5 gpc623_5_4787(
      {stage044[138], stage044[139], stage044[140]},
      {stage045[162], stage045[163]},
      {stage046[140], stage046[141], stage046[142], stage046[143], stage046[144], stage046[145]},
      {stage048[232], stage047[177], stage046[223], stage045[212], stage044[198]}
   );
   gpc623_5 gpc623_5_4788(
      {stage044[141], stage044[142], stage044[143]},
      {stage045[164], stage045[165]},
      {stage046[146], stage046[147], stage046[148], stage046[149], stage046[150], stage046[151]},
      {stage048[233], stage047[178], stage046[224], stage045[213], stage044[199]}
   );
   gpc623_5 gpc623_5_4789(
      {stage044[144], stage044[145], stage044[146]},
      {stage045[166], stage045[167]},
      {stage046[152], stage046[153], stage046[154], stage046[155], stage046[156], stage046[157]},
      {stage048[234], stage047[179], stage046[225], stage045[214], stage044[200]}
   );
   gpc623_5 gpc623_5_4790(
      {stage044[147], stage044[148], stage044[149]},
      {stage045[168], stage045[169]},
      {stage046[158], stage046[159], stage046[160], stage046[161], stage046[162], stage046[163]},
      {stage048[235], stage047[180], stage046[226], stage045[215], stage044[201]}
   );
   gpc623_5 gpc623_5_4791(
      {stage044[150], stage044[151], stage044[152]},
      {stage045[170], stage045[171]},
      {stage046[164], stage046[165], stage046[166], stage046[167], stage046[168], stage046[169]},
      {stage048[236], stage047[181], stage046[227], stage045[216], stage044[202]}
   );
   gpc606_5 gpc606_5_4792(
      {stage044[153], stage044[154], stage044[155], stage044[156], stage044[157], stage044[158]},
      {stage046[170], stage046[171], stage046[172], stage046[173], stage046[174], stage046[175]},
      {stage048[237], stage047[182], stage046[228], stage045[217], stage044[203]}
   );
   gpc615_5 gpc615_5_4793(
      {stage044[159], stage044[160], stage044[161], stage044[162], stage044[163]},
      {stage045[172]},
      {stage046[176], stage046[177], stage046[178], stage046[179], stage046[180], stage046[181]},
      {stage048[238], stage047[183], stage046[229], stage045[218], stage044[204]}
   );
   gpc615_5 gpc615_5_4794(
      {stage044[164], stage044[165], stage044[166], stage044[167], stage044[168]},
      {stage045[173]},
      {stage046[182], stage046[183], stage046[184], stage046[185], stage046[186], stage046[187]},
      {stage048[239], stage047[184], stage046[230], stage045[219], stage044[205]}
   );
   gpc615_5 gpc615_5_4795(
      {stage044[169], stage044[170], stage044[171], stage044[172], stage044[173]},
      {stage045[174]},
      {stage046[188], stage046[189], stage046[190], stage046[191], stage046[192], stage046[193]},
      {stage048[240], stage047[185], stage046[231], stage045[220], stage044[206]}
   );
   gpc615_5 gpc615_5_4796(
      {stage044[174], stage044[175], stage044[176], stage044[177], stage044[178]},
      {stage045[175]},
      {stage046[194], stage046[195], stage046[196], stage046[197], stage046[198], stage046[199]},
      {stage048[241], stage047[186], stage046[232], stage045[221], stage044[207]}
   );
   gpc1_1 gpc1_1_4797(
      {stage045[176]},
      {stage045[222]}
   );
   gpc1_1 gpc1_1_4798(
      {stage045[177]},
      {stage045[223]}
   );
   gpc1_1 gpc1_1_4799(
      {stage045[178]},
      {stage045[224]}
   );
   gpc1_1 gpc1_1_4800(
      {stage045[179]},
      {stage045[225]}
   );
   gpc1_1 gpc1_1_4801(
      {stage045[180]},
      {stage045[226]}
   );
   gpc1_1 gpc1_1_4802(
      {stage045[181]},
      {stage045[227]}
   );
   gpc1_1 gpc1_1_4803(
      {stage045[182]},
      {stage045[228]}
   );
   gpc1_1 gpc1_1_4804(
      {stage045[183]},
      {stage045[229]}
   );
   gpc1_1 gpc1_1_4805(
      {stage045[184]},
      {stage045[230]}
   );
   gpc1_1 gpc1_1_4806(
      {stage045[185]},
      {stage045[231]}
   );
   gpc1_1 gpc1_1_4807(
      {stage045[186]},
      {stage045[232]}
   );
   gpc1_1 gpc1_1_4808(
      {stage045[187]},
      {stage045[233]}
   );
   gpc1_1 gpc1_1_4809(
      {stage045[188]},
      {stage045[234]}
   );
   gpc1_1 gpc1_1_4810(
      {stage045[189]},
      {stage045[235]}
   );
   gpc1_1 gpc1_1_4811(
      {stage045[190]},
      {stage045[236]}
   );
   gpc1_1 gpc1_1_4812(
      {stage045[191]},
      {stage045[237]}
   );
   gpc1_1 gpc1_1_4813(
      {stage045[192]},
      {stage045[238]}
   );
   gpc1_1 gpc1_1_4814(
      {stage045[193]},
      {stage045[239]}
   );
   gpc1_1 gpc1_1_4815(
      {stage045[194]},
      {stage045[240]}
   );
   gpc1_1 gpc1_1_4816(
      {stage045[195]},
      {stage045[241]}
   );
   gpc1_1 gpc1_1_4817(
      {stage045[196]},
      {stage045[242]}
   );
   gpc1_1 gpc1_1_4818(
      {stage045[197]},
      {stage045[243]}
   );
   gpc1_1 gpc1_1_4819(
      {stage045[198]},
      {stage045[244]}
   );
   gpc1_1 gpc1_1_4820(
      {stage045[199]},
      {stage045[245]}
   );
   gpc1_1 gpc1_1_4821(
      {stage045[200]},
      {stage045[246]}
   );
   gpc1_1 gpc1_1_4822(
      {stage045[201]},
      {stage045[247]}
   );
   gpc1_1 gpc1_1_4823(
      {stage045[202]},
      {stage045[248]}
   );
   gpc1_1 gpc1_1_4824(
      {stage045[203]},
      {stage045[249]}
   );
   gpc1_1 gpc1_1_4825(
      {stage046[200]},
      {stage046[233]}
   );
   gpc1_1 gpc1_1_4826(
      {stage046[201]},
      {stage046[234]}
   );
   gpc1_1 gpc1_1_4827(
      {stage046[202]},
      {stage046[235]}
   );
   gpc1_1 gpc1_1_4828(
      {stage046[203]},
      {stage046[236]}
   );
   gpc1_1 gpc1_1_4829(
      {stage046[204]},
      {stage046[237]}
   );
   gpc1_1 gpc1_1_4830(
      {stage046[205]},
      {stage046[238]}
   );
   gpc1_1 gpc1_1_4831(
      {stage046[206]},
      {stage046[239]}
   );
   gpc1_1 gpc1_1_4832(
      {stage046[207]},
      {stage046[240]}
   );
   gpc1_1 gpc1_1_4833(
      {stage046[208]},
      {stage046[241]}
   );
   gpc1_1 gpc1_1_4834(
      {stage046[209]},
      {stage046[242]}
   );
   gpc1_1 gpc1_1_4835(
      {stage046[210]},
      {stage046[243]}
   );
   gpc1_1 gpc1_1_4836(
      {stage046[211]},
      {stage046[244]}
   );
   gpc1_1 gpc1_1_4837(
      {stage046[212]},
      {stage046[245]}
   );
   gpc1_1 gpc1_1_4838(
      {stage046[213]},
      {stage046[246]}
   );
   gpc1_1 gpc1_1_4839(
      {stage046[214]},
      {stage046[247]}
   );
   gpc1_1 gpc1_1_4840(
      {stage046[215]},
      {stage046[248]}
   );
   gpc623_5 gpc623_5_4841(
      {stage047[128], stage047[129], stage047[130]},
      {stage048[128], stage048[129]},
      {stage049[128], stage049[129], stage049[130], stage049[131], stage049[132], stage049[133]},
      {stage051[167], stage050[224], stage049[204], stage048[242], stage047[187]}
   );
   gpc623_5 gpc623_5_4842(
      {stage047[131], stage047[132], stage047[133]},
      {stage048[130], stage048[131]},
      {stage049[134], stage049[135], stage049[136], stage049[137], stage049[138], stage049[139]},
      {stage051[168], stage050[225], stage049[205], stage048[243], stage047[188]}
   );
   gpc623_5 gpc623_5_4843(
      {stage047[134], stage047[135], stage047[136]},
      {stage048[132], stage048[133]},
      {stage049[140], stage049[141], stage049[142], stage049[143], stage049[144], stage049[145]},
      {stage051[169], stage050[226], stage049[206], stage048[244], stage047[189]}
   );
   gpc623_5 gpc623_5_4844(
      {stage047[137], stage047[138], stage047[139]},
      {stage048[134], stage048[135]},
      {stage049[146], stage049[147], stage049[148], stage049[149], stage049[150], stage049[151]},
      {stage051[170], stage050[227], stage049[207], stage048[245], stage047[190]}
   );
   gpc623_5 gpc623_5_4845(
      {stage047[140], stage047[141], stage047[142]},
      {stage048[136], stage048[137]},
      {stage049[152], stage049[153], stage049[154], stage049[155], stage049[156], stage049[157]},
      {stage051[171], stage050[228], stage049[208], stage048[246], stage047[191]}
   );
   gpc623_5 gpc623_5_4846(
      {stage047[143], stage047[144], stage047[145]},
      {stage048[138], stage048[139]},
      {stage049[158], stage049[159], stage049[160], stage049[161], stage049[162], stage049[163]},
      {stage051[172], stage050[229], stage049[209], stage048[247], stage047[192]}
   );
   gpc615_5 gpc615_5_4847(
      {stage047[146], stage047[147], stage047[148], stage047[149], stage047[150]},
      {stage048[140]},
      {stage049[164], stage049[165], stage049[166], stage049[167], stage049[168], stage049[169]},
      {stage051[173], stage050[230], stage049[210], stage048[248], stage047[193]}
   );
   gpc615_5 gpc615_5_4848(
      {stage047[151], stage047[152], stage047[153], stage047[154], stage047[155]},
      {stage048[141]},
      {stage049[170], stage049[171], stage049[172], stage049[173], stage049[174], stage049[175]},
      {stage051[174], stage050[231], stage049[211], stage048[249], stage047[194]}
   );
   gpc615_5 gpc615_5_4849(
      {stage047[156], stage047[157], stage047[158], stage047[159], stage047[160]},
      {stage048[142]},
      {stage049[176], stage049[177], stage049[178], stage049[179], stage049[180], stage049[181]},
      {stage051[175], stage050[232], stage049[212], stage048[250], stage047[195]}
   );
   gpc615_5 gpc615_5_4850(
      {stage047[161], stage047[162], stage047[163], stage047[164], stage047[165]},
      {stage048[143]},
      {stage049[182], stage049[183], stage049[184], stage049[185], stage049[186], stage049[187]},
      {stage051[176], stage050[233], stage049[213], stage048[251], stage047[196]}
   );
   gpc615_5 gpc615_5_4851(
      {stage047[166], stage047[167], stage047[168], stage047[169], 1'h0},
      {stage048[144]},
      {stage049[188], stage049[189], stage049[190], stage049[191], stage049[192], stage049[193]},
      {stage051[177], stage050[234], stage049[214], stage048[252], stage047[197]}
   );
   gpc1_1 gpc1_1_4852(
      {stage048[145]},
      {stage048[253]}
   );
   gpc1_1 gpc1_1_4853(
      {stage048[146]},
      {stage048[254]}
   );
   gpc1_1 gpc1_1_4854(
      {stage048[147]},
      {stage048[255]}
   );
   gpc1_1 gpc1_1_4855(
      {stage048[148]},
      {stage048[256]}
   );
   gpc1_1 gpc1_1_4856(
      {stage048[149]},
      {stage048[257]}
   );
   gpc1_1 gpc1_1_4857(
      {stage048[150]},
      {stage048[258]}
   );
   gpc1_1 gpc1_1_4858(
      {stage048[151]},
      {stage048[259]}
   );
   gpc1_1 gpc1_1_4859(
      {stage048[152]},
      {stage048[260]}
   );
   gpc1_1 gpc1_1_4860(
      {stage048[153]},
      {stage048[261]}
   );
   gpc1_1 gpc1_1_4861(
      {stage048[154]},
      {stage048[262]}
   );
   gpc1_1 gpc1_1_4862(
      {stage048[155]},
      {stage048[263]}
   );
   gpc1_1 gpc1_1_4863(
      {stage048[156]},
      {stage048[264]}
   );
   gpc1_1 gpc1_1_4864(
      {stage048[157]},
      {stage048[265]}
   );
   gpc1_1 gpc1_1_4865(
      {stage048[158]},
      {stage048[266]}
   );
   gpc1_1 gpc1_1_4866(
      {stage048[159]},
      {stage048[267]}
   );
   gpc1_1 gpc1_1_4867(
      {stage048[160]},
      {stage048[268]}
   );
   gpc1_1 gpc1_1_4868(
      {stage048[161]},
      {stage048[269]}
   );
   gpc1_1 gpc1_1_4869(
      {stage048[162]},
      {stage048[270]}
   );
   gpc1_1 gpc1_1_4870(
      {stage048[163]},
      {stage048[271]}
   );
   gpc1_1 gpc1_1_4871(
      {stage048[164]},
      {stage048[272]}
   );
   gpc1_1 gpc1_1_4872(
      {stage048[165]},
      {stage048[273]}
   );
   gpc1_1 gpc1_1_4873(
      {stage048[166]},
      {stage048[274]}
   );
   gpc1_1 gpc1_1_4874(
      {stage048[167]},
      {stage048[275]}
   );
   gpc1_1 gpc1_1_4875(
      {stage048[168]},
      {stage048[276]}
   );
   gpc1_1 gpc1_1_4876(
      {stage048[169]},
      {stage048[277]}
   );
   gpc1_1 gpc1_1_4877(
      {stage048[170]},
      {stage048[278]}
   );
   gpc1_1 gpc1_1_4878(
      {stage048[171]},
      {stage048[279]}
   );
   gpc1_1 gpc1_1_4879(
      {stage048[172]},
      {stage048[280]}
   );
   gpc1_1 gpc1_1_4880(
      {stage048[173]},
      {stage048[281]}
   );
   gpc1_1 gpc1_1_4881(
      {stage048[174]},
      {stage048[282]}
   );
   gpc1_1 gpc1_1_4882(
      {stage048[175]},
      {stage048[283]}
   );
   gpc1_1 gpc1_1_4883(
      {stage048[176]},
      {stage048[284]}
   );
   gpc1_1 gpc1_1_4884(
      {stage048[177]},
      {stage048[285]}
   );
   gpc606_5 gpc606_5_4885(
      {stage048[178], stage048[179], stage048[180], stage048[181], stage048[182], stage048[183]},
      {stage050[128], stage050[129], stage050[130], stage050[131], stage050[132], stage050[133]},
      {stage052[214], stage051[178], stage050[235], stage049[215], stage048[286]}
   );
   gpc606_5 gpc606_5_4886(
      {stage048[184], stage048[185], stage048[186], stage048[187], stage048[188], stage048[189]},
      {stage050[134], stage050[135], stage050[136], stage050[137], stage050[138], stage050[139]},
      {stage052[215], stage051[179], stage050[236], stage049[216], stage048[287]}
   );
   gpc606_5 gpc606_5_4887(
      {stage048[190], stage048[191], stage048[192], stage048[193], stage048[194], stage048[195]},
      {stage050[140], stage050[141], stage050[142], stage050[143], stage050[144], stage050[145]},
      {stage052[216], stage051[180], stage050[237], stage049[217], stage048[288]}
   );
   gpc606_5 gpc606_5_4888(
      {stage048[196], stage048[197], stage048[198], stage048[199], stage048[200], stage048[201]},
      {stage050[146], stage050[147], stage050[148], stage050[149], stage050[150], stage050[151]},
      {stage052[217], stage051[181], stage050[238], stage049[218], stage048[289]}
   );
   gpc606_5 gpc606_5_4889(
      {stage048[202], stage048[203], stage048[204], stage048[205], stage048[206], stage048[207]},
      {stage050[152], stage050[153], stage050[154], stage050[155], stage050[156], stage050[157]},
      {stage052[218], stage051[182], stage050[239], stage049[219], stage048[290]}
   );
   gpc606_5 gpc606_5_4890(
      {stage048[208], stage048[209], stage048[210], stage048[211], stage048[212], stage048[213]},
      {stage050[158], stage050[159], stage050[160], stage050[161], stage050[162], stage050[163]},
      {stage052[219], stage051[183], stage050[240], stage049[220], stage048[291]}
   );
   gpc606_5 gpc606_5_4891(
      {stage048[214], stage048[215], stage048[216], stage048[217], stage048[218], stage048[219]},
      {stage050[164], stage050[165], stage050[166], stage050[167], stage050[168], stage050[169]},
      {stage052[220], stage051[184], stage050[241], stage049[221], stage048[292]}
   );
   gpc615_5 gpc615_5_4892(
      {stage048[220], stage048[221], stage048[222], stage048[223], stage048[224]},
      {stage049[194]},
      {stage050[170], stage050[171], stage050[172], stage050[173], stage050[174], stage050[175]},
      {stage052[221], stage051[185], stage050[242], stage049[222], stage048[293]}
   );
   gpc135_4 gpc135_4_4893(
      {stage048[225], stage048[226], stage048[227], stage048[228], stage048[229]},
      {stage049[195], stage049[196], stage049[197]},
      {stage050[176]},
      {stage051[186], stage050[243], stage049[223], stage048[294]}
   );
   gpc1_1 gpc1_1_4894(
      {stage049[198]},
      {stage049[224]}
   );
   gpc1_1 gpc1_1_4895(
      {stage049[199]},
      {stage049[225]}
   );
   gpc1_1 gpc1_1_4896(
      {stage049[200]},
      {stage049[226]}
   );
   gpc1_1 gpc1_1_4897(
      {stage049[201]},
      {stage049[227]}
   );
   gpc1_1 gpc1_1_4898(
      {stage049[202]},
      {stage049[228]}
   );
   gpc1_1 gpc1_1_4899(
      {stage049[203]},
      {stage049[229]}
   );
   gpc1_1 gpc1_1_4900(
      {stage050[177]},
      {stage050[244]}
   );
   gpc1_1 gpc1_1_4901(
      {stage050[178]},
      {stage050[245]}
   );
   gpc615_5 gpc615_5_4902(
      {stage050[179], stage050[180], stage050[181], stage050[182], stage050[183]},
      {stage051[128]},
      {stage052[128], stage052[129], stage052[130], stage052[131], stage052[132], stage052[133]},
      {stage054[205], stage053[171], stage052[222], stage051[187], stage050[246]}
   );
   gpc615_5 gpc615_5_4903(
      {stage050[184], stage050[185], stage050[186], stage050[187], stage050[188]},
      {stage051[129]},
      {stage052[134], stage052[135], stage052[136], stage052[137], stage052[138], stage052[139]},
      {stage054[206], stage053[172], stage052[223], stage051[188], stage050[247]}
   );
   gpc615_5 gpc615_5_4904(
      {stage050[189], stage050[190], stage050[191], stage050[192], stage050[193]},
      {stage051[130]},
      {stage052[140], stage052[141], stage052[142], stage052[143], stage052[144], stage052[145]},
      {stage054[207], stage053[173], stage052[224], stage051[189], stage050[248]}
   );
   gpc615_5 gpc615_5_4905(
      {stage050[194], stage050[195], stage050[196], stage050[197], stage050[198]},
      {stage051[131]},
      {stage052[146], stage052[147], stage052[148], stage052[149], stage052[150], stage052[151]},
      {stage054[208], stage053[174], stage052[225], stage051[190], stage050[249]}
   );
   gpc615_5 gpc615_5_4906(
      {stage050[199], stage050[200], stage050[201], stage050[202], stage050[203]},
      {stage051[132]},
      {stage052[152], stage052[153], stage052[154], stage052[155], stage052[156], stage052[157]},
      {stage054[209], stage053[175], stage052[226], stage051[191], stage050[250]}
   );
   gpc615_5 gpc615_5_4907(
      {stage050[204], stage050[205], stage050[206], stage050[207], stage050[208]},
      {stage051[133]},
      {stage052[158], stage052[159], stage052[160], stage052[161], stage052[162], stage052[163]},
      {stage054[210], stage053[176], stage052[227], stage051[192], stage050[251]}
   );
   gpc615_5 gpc615_5_4908(
      {stage050[209], stage050[210], stage050[211], stage050[212], stage050[213]},
      {stage051[134]},
      {stage052[164], stage052[165], stage052[166], stage052[167], stage052[168], stage052[169]},
      {stage054[211], stage053[177], stage052[228], stage051[193], stage050[252]}
   );
   gpc615_5 gpc615_5_4909(
      {stage050[214], stage050[215], stage050[216], stage050[217], stage050[218]},
      {stage051[135]},
      {stage052[170], stage052[171], stage052[172], stage052[173], stage052[174], stage052[175]},
      {stage054[212], stage053[178], stage052[229], stage051[194], stage050[253]}
   );
   gpc615_5 gpc615_5_4910(
      {stage050[219], stage050[220], stage050[221], stage050[222], stage050[223]},
      {stage051[136]},
      {stage052[176], stage052[177], stage052[178], stage052[179], stage052[180], stage052[181]},
      {stage054[213], stage053[179], stage052[230], stage051[195], stage050[254]}
   );
   gpc1_1 gpc1_1_4911(
      {stage051[137]},
      {stage051[196]}
   );
   gpc1_1 gpc1_1_4912(
      {stage051[138]},
      {stage051[197]}
   );
   gpc1_1 gpc1_1_4913(
      {stage051[139]},
      {stage051[198]}
   );
   gpc1_1 gpc1_1_4914(
      {stage051[140]},
      {stage051[199]}
   );
   gpc1_1 gpc1_1_4915(
      {stage051[141]},
      {stage051[200]}
   );
   gpc1_1 gpc1_1_4916(
      {stage051[142]},
      {stage051[201]}
   );
   gpc1_1 gpc1_1_4917(
      {stage051[143]},
      {stage051[202]}
   );
   gpc1_1 gpc1_1_4918(
      {stage051[144]},
      {stage051[203]}
   );
   gpc1_1 gpc1_1_4919(
      {stage051[145]},
      {stage051[204]}
   );
   gpc1_1 gpc1_1_4920(
      {stage051[146]},
      {stage051[205]}
   );
   gpc1_1 gpc1_1_4921(
      {stage051[147]},
      {stage051[206]}
   );
   gpc1_1 gpc1_1_4922(
      {stage051[148]},
      {stage051[207]}
   );
   gpc1_1 gpc1_1_4923(
      {stage051[149]},
      {stage051[208]}
   );
   gpc1_1 gpc1_1_4924(
      {stage051[150]},
      {stage051[209]}
   );
   gpc1_1 gpc1_1_4925(
      {stage051[151]},
      {stage051[210]}
   );
   gpc1_1 gpc1_1_4926(
      {stage051[152]},
      {stage051[211]}
   );
   gpc1_1 gpc1_1_4927(
      {stage051[153]},
      {stage051[212]}
   );
   gpc1_1 gpc1_1_4928(
      {stage051[154]},
      {stage051[213]}
   );
   gpc1_1 gpc1_1_4929(
      {stage051[155]},
      {stage051[214]}
   );
   gpc1_1 gpc1_1_4930(
      {stage051[156]},
      {stage051[215]}
   );
   gpc1_1 gpc1_1_4931(
      {stage051[157]},
      {stage051[216]}
   );
   gpc1_1 gpc1_1_4932(
      {stage051[158]},
      {stage051[217]}
   );
   gpc1_1 gpc1_1_4933(
      {stage051[159]},
      {stage051[218]}
   );
   gpc1_1 gpc1_1_4934(
      {stage051[160]},
      {stage051[219]}
   );
   gpc1_1 gpc1_1_4935(
      {stage051[161]},
      {stage051[220]}
   );
   gpc615_5 gpc615_5_4936(
      {stage051[162], stage051[163], stage051[164], stage051[165], stage051[166]},
      {stage052[182]},
      {stage053[128], stage053[129], stage053[130], stage053[131], stage053[132], stage053[133]},
      {stage055[199], stage054[214], stage053[180], stage052[231], stage051[221]}
   );
   gpc1_1 gpc1_1_4937(
      {stage052[183]},
      {stage052[232]}
   );
   gpc1_1 gpc1_1_4938(
      {stage052[184]},
      {stage052[233]}
   );
   gpc1_1 gpc1_1_4939(
      {stage052[185]},
      {stage052[234]}
   );
   gpc1_1 gpc1_1_4940(
      {stage052[186]},
      {stage052[235]}
   );
   gpc1_1 gpc1_1_4941(
      {stage052[187]},
      {stage052[236]}
   );
   gpc1_1 gpc1_1_4942(
      {stage052[188]},
      {stage052[237]}
   );
   gpc1_1 gpc1_1_4943(
      {stage052[189]},
      {stage052[238]}
   );
   gpc606_5 gpc606_5_4944(
      {stage052[190], stage052[191], stage052[192], stage052[193], stage052[194], stage052[195]},
      {stage054[128], stage054[129], stage054[130], stage054[131], stage054[132], stage054[133]},
      {stage056[205], stage055[200], stage054[215], stage053[181], stage052[239]}
   );
   gpc606_5 gpc606_5_4945(
      {stage052[196], stage052[197], stage052[198], stage052[199], stage052[200], stage052[201]},
      {stage054[134], stage054[135], stage054[136], stage054[137], stage054[138], stage054[139]},
      {stage056[206], stage055[201], stage054[216], stage053[182], stage052[240]}
   );
   gpc606_5 gpc606_5_4946(
      {stage052[202], stage052[203], stage052[204], stage052[205], stage052[206], stage052[207]},
      {stage054[140], stage054[141], stage054[142], stage054[143], stage054[144], stage054[145]},
      {stage056[207], stage055[202], stage054[217], stage053[183], stage052[241]}
   );
   gpc606_5 gpc606_5_4947(
      {stage052[208], stage052[209], stage052[210], stage052[211], stage052[212], stage052[213]},
      {stage054[146], stage054[147], stage054[148], stage054[149], stage054[150], stage054[151]},
      {stage056[208], stage055[203], stage054[218], stage053[184], stage052[242]}
   );
   gpc1_1 gpc1_1_4948(
      {stage053[134]},
      {stage053[185]}
   );
   gpc1_1 gpc1_1_4949(
      {stage053[135]},
      {stage053[186]}
   );
   gpc1_1 gpc1_1_4950(
      {stage053[136]},
      {stage053[187]}
   );
   gpc1_1 gpc1_1_4951(
      {stage053[137]},
      {stage053[188]}
   );
   gpc1_1 gpc1_1_4952(
      {stage053[138]},
      {stage053[189]}
   );
   gpc1_1 gpc1_1_4953(
      {stage053[139]},
      {stage053[190]}
   );
   gpc1_1 gpc1_1_4954(
      {stage053[140]},
      {stage053[191]}
   );
   gpc1_1 gpc1_1_4955(
      {stage053[141]},
      {stage053[192]}
   );
   gpc1_1 gpc1_1_4956(
      {stage053[142]},
      {stage053[193]}
   );
   gpc1_1 gpc1_1_4957(
      {stage053[143]},
      {stage053[194]}
   );
   gpc1_1 gpc1_1_4958(
      {stage053[144]},
      {stage053[195]}
   );
   gpc1_1 gpc1_1_4959(
      {stage053[145]},
      {stage053[196]}
   );
   gpc1_1 gpc1_1_4960(
      {stage053[146]},
      {stage053[197]}
   );
   gpc1_1 gpc1_1_4961(
      {stage053[147]},
      {stage053[198]}
   );
   gpc1_1 gpc1_1_4962(
      {stage053[148]},
      {stage053[199]}
   );
   gpc1_1 gpc1_1_4963(
      {stage053[149]},
      {stage053[200]}
   );
   gpc1_1 gpc1_1_4964(
      {stage053[150]},
      {stage053[201]}
   );
   gpc1_1 gpc1_1_4965(
      {stage053[151]},
      {stage053[202]}
   );
   gpc1_1 gpc1_1_4966(
      {stage053[152]},
      {stage053[203]}
   );
   gpc1_1 gpc1_1_4967(
      {stage053[153]},
      {stage053[204]}
   );
   gpc1_1 gpc1_1_4968(
      {stage053[154]},
      {stage053[205]}
   );
   gpc1_1 gpc1_1_4969(
      {stage053[155]},
      {stage053[206]}
   );
   gpc1_1 gpc1_1_4970(
      {stage053[156]},
      {stage053[207]}
   );
   gpc1_1 gpc1_1_4971(
      {stage053[157]},
      {stage053[208]}
   );
   gpc1_1 gpc1_1_4972(
      {stage053[158]},
      {stage053[209]}
   );
   gpc606_5 gpc606_5_4973(
      {stage053[159], stage053[160], stage053[161], stage053[162], stage053[163], stage053[164]},
      {stage055[128], stage055[129], stage055[130], stage055[131], stage055[132], stage055[133]},
      {stage057[184], stage056[209], stage055[204], stage054[219], stage053[210]}
   );
   gpc606_5 gpc606_5_4974(
      {stage053[165], stage053[166], stage053[167], stage053[168], stage053[169], stage053[170]},
      {stage055[134], stage055[135], stage055[136], stage055[137], stage055[138], stage055[139]},
      {stage057[185], stage056[210], stage055[205], stage054[220], stage053[211]}
   );
   gpc1_1 gpc1_1_4975(
      {stage054[152]},
      {stage054[221]}
   );
   gpc1_1 gpc1_1_4976(
      {stage054[153]},
      {stage054[222]}
   );
   gpc1_1 gpc1_1_4977(
      {stage054[154]},
      {stage054[223]}
   );
   gpc615_5 gpc615_5_4978(
      {stage054[155], stage054[156], stage054[157], stage054[158], stage054[159]},
      {stage055[140]},
      {stage056[128], stage056[129], stage056[130], stage056[131], stage056[132], stage056[133]},
      {stage058[180], stage057[186], stage056[211], stage055[206], stage054[224]}
   );
   gpc615_5 gpc615_5_4979(
      {stage054[160], stage054[161], stage054[162], stage054[163], stage054[164]},
      {stage055[141]},
      {stage056[134], stage056[135], stage056[136], stage056[137], stage056[138], stage056[139]},
      {stage058[181], stage057[187], stage056[212], stage055[207], stage054[225]}
   );
   gpc615_5 gpc615_5_4980(
      {stage054[165], stage054[166], stage054[167], stage054[168], stage054[169]},
      {stage055[142]},
      {stage056[140], stage056[141], stage056[142], stage056[143], stage056[144], stage056[145]},
      {stage058[182], stage057[188], stage056[213], stage055[208], stage054[226]}
   );
   gpc615_5 gpc615_5_4981(
      {stage054[170], stage054[171], stage054[172], stage054[173], stage054[174]},
      {stage055[143]},
      {stage056[146], stage056[147], stage056[148], stage056[149], stage056[150], stage056[151]},
      {stage058[183], stage057[189], stage056[214], stage055[209], stage054[227]}
   );
   gpc615_5 gpc615_5_4982(
      {stage054[175], stage054[176], stage054[177], stage054[178], stage054[179]},
      {stage055[144]},
      {stage056[152], stage056[153], stage056[154], stage056[155], stage056[156], stage056[157]},
      {stage058[184], stage057[190], stage056[215], stage055[210], stage054[228]}
   );
   gpc615_5 gpc615_5_4983(
      {stage054[180], stage054[181], stage054[182], stage054[183], stage054[184]},
      {stage055[145]},
      {stage056[158], stage056[159], stage056[160], stage056[161], stage056[162], stage056[163]},
      {stage058[185], stage057[191], stage056[216], stage055[211], stage054[229]}
   );
   gpc615_5 gpc615_5_4984(
      {stage054[185], stage054[186], stage054[187], stage054[188], stage054[189]},
      {stage055[146]},
      {stage056[164], stage056[165], stage056[166], stage056[167], stage056[168], stage056[169]},
      {stage058[186], stage057[192], stage056[217], stage055[212], stage054[230]}
   );
   gpc615_5 gpc615_5_4985(
      {stage054[190], stage054[191], stage054[192], stage054[193], stage054[194]},
      {stage055[147]},
      {stage056[170], stage056[171], stage056[172], stage056[173], stage056[174], stage056[175]},
      {stage058[187], stage057[193], stage056[218], stage055[213], stage054[231]}
   );
   gpc615_5 gpc615_5_4986(
      {stage054[195], stage054[196], stage054[197], stage054[198], stage054[199]},
      {stage055[148]},
      {stage056[176], stage056[177], stage056[178], stage056[179], stage056[180], stage056[181]},
      {stage058[188], stage057[194], stage056[219], stage055[214], stage054[232]}
   );
   gpc615_5 gpc615_5_4987(
      {stage054[200], stage054[201], stage054[202], stage054[203], stage054[204]},
      {stage055[149]},
      {stage056[182], stage056[183], stage056[184], stage056[185], stage056[186], stage056[187]},
      {stage058[189], stage057[195], stage056[220], stage055[215], stage054[233]}
   );
   gpc1_1 gpc1_1_4988(
      {stage055[150]},
      {stage055[216]}
   );
   gpc1_1 gpc1_1_4989(
      {stage055[151]},
      {stage055[217]}
   );
   gpc1_1 gpc1_1_4990(
      {stage055[152]},
      {stage055[218]}
   );
   gpc1_1 gpc1_1_4991(
      {stage055[153]},
      {stage055[219]}
   );
   gpc1_1 gpc1_1_4992(
      {stage055[154]},
      {stage055[220]}
   );
   gpc1_1 gpc1_1_4993(
      {stage055[155]},
      {stage055[221]}
   );
   gpc1_1 gpc1_1_4994(
      {stage055[156]},
      {stage055[222]}
   );
   gpc1_1 gpc1_1_4995(
      {stage055[157]},
      {stage055[223]}
   );
   gpc1_1 gpc1_1_4996(
      {stage055[158]},
      {stage055[224]}
   );
   gpc1_1 gpc1_1_4997(
      {stage055[159]},
      {stage055[225]}
   );
   gpc1_1 gpc1_1_4998(
      {stage055[160]},
      {stage055[226]}
   );
   gpc1_1 gpc1_1_4999(
      {stage055[161]},
      {stage055[227]}
   );
   gpc1_1 gpc1_1_5000(
      {stage055[162]},
      {stage055[228]}
   );
   gpc1_1 gpc1_1_5001(
      {stage055[163]},
      {stage055[229]}
   );
   gpc1_1 gpc1_1_5002(
      {stage055[164]},
      {stage055[230]}
   );
   gpc1_1 gpc1_1_5003(
      {stage055[165]},
      {stage055[231]}
   );
   gpc1_1 gpc1_1_5004(
      {stage055[166]},
      {stage055[232]}
   );
   gpc1_1 gpc1_1_5005(
      {stage055[167]},
      {stage055[233]}
   );
   gpc1_1 gpc1_1_5006(
      {stage055[168]},
      {stage055[234]}
   );
   gpc1_1 gpc1_1_5007(
      {stage055[169]},
      {stage055[235]}
   );
   gpc1_1 gpc1_1_5008(
      {stage055[170]},
      {stage055[236]}
   );
   gpc1_1 gpc1_1_5009(
      {stage055[171]},
      {stage055[237]}
   );
   gpc1_1 gpc1_1_5010(
      {stage055[172]},
      {stage055[238]}
   );
   gpc1_1 gpc1_1_5011(
      {stage055[173]},
      {stage055[239]}
   );
   gpc1_1 gpc1_1_5012(
      {stage055[174]},
      {stage055[240]}
   );
   gpc1_1 gpc1_1_5013(
      {stage055[175]},
      {stage055[241]}
   );
   gpc1_1 gpc1_1_5014(
      {stage055[176]},
      {stage055[242]}
   );
   gpc606_5 gpc606_5_5015(
      {stage055[177], stage055[178], stage055[179], stage055[180], stage055[181], stage055[182]},
      {stage057[128], stage057[129], stage057[130], stage057[131], stage057[132], stage057[133]},
      {stage059[216], stage058[190], stage057[196], stage056[221], stage055[243]}
   );
   gpc606_5 gpc606_5_5016(
      {stage055[183], stage055[184], stage055[185], stage055[186], stage055[187], stage055[188]},
      {stage057[134], stage057[135], stage057[136], stage057[137], stage057[138], stage057[139]},
      {stage059[217], stage058[191], stage057[197], stage056[222], stage055[244]}
   );
   gpc615_5 gpc615_5_5017(
      {stage055[189], stage055[190], stage055[191], stage055[192], stage055[193]},
      {stage056[188]},
      {stage057[140], stage057[141], stage057[142], stage057[143], stage057[144], stage057[145]},
      {stage059[218], stage058[192], stage057[198], stage056[223], stage055[245]}
   );
   gpc615_5 gpc615_5_5018(
      {stage055[194], stage055[195], stage055[196], stage055[197], stage055[198]},
      {stage056[189]},
      {stage057[146], stage057[147], stage057[148], stage057[149], stage057[150], stage057[151]},
      {stage059[219], stage058[193], stage057[199], stage056[224], stage055[246]}
   );
   gpc1_1 gpc1_1_5019(
      {stage056[190]},
      {stage056[225]}
   );
   gpc1_1 gpc1_1_5020(
      {stage056[191]},
      {stage056[226]}
   );
   gpc1_1 gpc1_1_5021(
      {stage056[192]},
      {stage056[227]}
   );
   gpc1_1 gpc1_1_5022(
      {stage056[193]},
      {stage056[228]}
   );
   gpc1_1 gpc1_1_5023(
      {stage056[194]},
      {stage056[229]}
   );
   gpc1_1 gpc1_1_5024(
      {stage056[195]},
      {stage056[230]}
   );
   gpc1_1 gpc1_1_5025(
      {stage056[196]},
      {stage056[231]}
   );
   gpc1_1 gpc1_1_5026(
      {stage056[197]},
      {stage056[232]}
   );
   gpc1_1 gpc1_1_5027(
      {stage056[198]},
      {stage056[233]}
   );
   gpc606_5 gpc606_5_5028(
      {stage056[199], stage056[200], stage056[201], stage056[202], stage056[203], stage056[204]},
      {stage058[128], stage058[129], stage058[130], stage058[131], stage058[132], stage058[133]},
      {stage060[190], stage059[220], stage058[194], stage057[200], stage056[234]}
   );
   gpc1_1 gpc1_1_5029(
      {stage057[152]},
      {stage057[201]}
   );
   gpc1_1 gpc1_1_5030(
      {stage057[153]},
      {stage057[202]}
   );
   gpc1_1 gpc1_1_5031(
      {stage057[154]},
      {stage057[203]}
   );
   gpc1_1 gpc1_1_5032(
      {stage057[155]},
      {stage057[204]}
   );
   gpc1_1 gpc1_1_5033(
      {stage057[156]},
      {stage057[205]}
   );
   gpc1_1 gpc1_1_5034(
      {stage057[157]},
      {stage057[206]}
   );
   gpc1_1 gpc1_1_5035(
      {stage057[158]},
      {stage057[207]}
   );
   gpc1_1 gpc1_1_5036(
      {stage057[159]},
      {stage057[208]}
   );
   gpc1_1 gpc1_1_5037(
      {stage057[160]},
      {stage057[209]}
   );
   gpc1_1 gpc1_1_5038(
      {stage057[161]},
      {stage057[210]}
   );
   gpc1_1 gpc1_1_5039(
      {stage057[162]},
      {stage057[211]}
   );
   gpc1_1 gpc1_1_5040(
      {stage057[163]},
      {stage057[212]}
   );
   gpc1_1 gpc1_1_5041(
      {stage057[164]},
      {stage057[213]}
   );
   gpc1_1 gpc1_1_5042(
      {stage057[165]},
      {stage057[214]}
   );
   gpc1_1 gpc1_1_5043(
      {stage057[166]},
      {stage057[215]}
   );
   gpc1_1 gpc1_1_5044(
      {stage057[167]},
      {stage057[216]}
   );
   gpc1_1 gpc1_1_5045(
      {stage057[168]},
      {stage057[217]}
   );
   gpc1_1 gpc1_1_5046(
      {stage057[169]},
      {stage057[218]}
   );
   gpc1_1 gpc1_1_5047(
      {stage057[170]},
      {stage057[219]}
   );
   gpc1_1 gpc1_1_5048(
      {stage057[171]},
      {stage057[220]}
   );
   gpc1_1 gpc1_1_5049(
      {stage057[172]},
      {stage057[221]}
   );
   gpc1_1 gpc1_1_5050(
      {stage057[173]},
      {stage057[222]}
   );
   gpc1_1 gpc1_1_5051(
      {stage057[174]},
      {stage057[223]}
   );
   gpc1_1 gpc1_1_5052(
      {stage057[175]},
      {stage057[224]}
   );
   gpc1_1 gpc1_1_5053(
      {stage057[176]},
      {stage057[225]}
   );
   gpc1_1 gpc1_1_5054(
      {stage057[177]},
      {stage057[226]}
   );
   gpc1_1 gpc1_1_5055(
      {stage057[178]},
      {stage057[227]}
   );
   gpc1_1 gpc1_1_5056(
      {stage057[179]},
      {stage057[228]}
   );
   gpc1_1 gpc1_1_5057(
      {stage057[180]},
      {stage057[229]}
   );
   gpc1_1 gpc1_1_5058(
      {stage057[181]},
      {stage057[230]}
   );
   gpc1_1 gpc1_1_5059(
      {stage057[182]},
      {stage057[231]}
   );
   gpc1_1 gpc1_1_5060(
      {stage057[183]},
      {stage057[232]}
   );
   gpc1_1 gpc1_1_5061(
      {stage058[134]},
      {stage058[195]}
   );
   gpc1_1 gpc1_1_5062(
      {stage058[135]},
      {stage058[196]}
   );
   gpc1_1 gpc1_1_5063(
      {stage058[136]},
      {stage058[197]}
   );
   gpc1_1 gpc1_1_5064(
      {stage058[137]},
      {stage058[198]}
   );
   gpc1_1 gpc1_1_5065(
      {stage058[138]},
      {stage058[199]}
   );
   gpc1_1 gpc1_1_5066(
      {stage058[139]},
      {stage058[200]}
   );
   gpc615_5 gpc615_5_5067(
      {stage058[140], stage058[141], stage058[142], stage058[143], stage058[144]},
      {stage059[128]},
      {stage060[128], stage060[129], stage060[130], stage060[131], stage060[132], stage060[133]},
      {stage062[189], stage061[189], stage060[191], stage059[221], stage058[201]}
   );
   gpc615_5 gpc615_5_5068(
      {stage058[145], stage058[146], stage058[147], stage058[148], stage058[149]},
      {stage059[129]},
      {stage060[134], stage060[135], stage060[136], stage060[137], stage060[138], stage060[139]},
      {stage062[190], stage061[190], stage060[192], stage059[222], stage058[202]}
   );
   gpc615_5 gpc615_5_5069(
      {stage058[150], stage058[151], stage058[152], stage058[153], stage058[154]},
      {stage059[130]},
      {stage060[140], stage060[141], stage060[142], stage060[143], stage060[144], stage060[145]},
      {stage062[191], stage061[191], stage060[193], stage059[223], stage058[203]}
   );
   gpc615_5 gpc615_5_5070(
      {stage058[155], stage058[156], stage058[157], stage058[158], stage058[159]},
      {stage059[131]},
      {stage060[146], stage060[147], stage060[148], stage060[149], stage060[150], stage060[151]},
      {stage062[192], stage061[192], stage060[194], stage059[224], stage058[204]}
   );
   gpc615_5 gpc615_5_5071(
      {stage058[160], stage058[161], stage058[162], stage058[163], stage058[164]},
      {stage059[132]},
      {stage060[152], stage060[153], stage060[154], stage060[155], stage060[156], stage060[157]},
      {stage062[193], stage061[193], stage060[195], stage059[225], stage058[205]}
   );
   gpc615_5 gpc615_5_5072(
      {stage058[165], stage058[166], stage058[167], stage058[168], stage058[169]},
      {stage059[133]},
      {stage060[158], stage060[159], stage060[160], stage060[161], stage060[162], stage060[163]},
      {stage062[194], stage061[194], stage060[196], stage059[226], stage058[206]}
   );
   gpc615_5 gpc615_5_5073(
      {stage058[170], stage058[171], stage058[172], stage058[173], stage058[174]},
      {stage059[134]},
      {stage060[164], stage060[165], stage060[166], stage060[167], stage060[168], stage060[169]},
      {stage062[195], stage061[195], stage060[197], stage059[227], stage058[207]}
   );
   gpc615_5 gpc615_5_5074(
      {stage058[175], stage058[176], stage058[177], stage058[178], stage058[179]},
      {stage059[135]},
      {stage060[170], stage060[171], stage060[172], stage060[173], stage060[174], stage060[175]},
      {stage062[196], stage061[196], stage060[198], stage059[228], stage058[208]}
   );
   gpc1_1 gpc1_1_5075(
      {stage059[136]},
      {stage059[229]}
   );
   gpc1_1 gpc1_1_5076(
      {stage059[137]},
      {stage059[230]}
   );
   gpc1_1 gpc1_1_5077(
      {stage059[138]},
      {stage059[231]}
   );
   gpc1_1 gpc1_1_5078(
      {stage059[139]},
      {stage059[232]}
   );
   gpc1_1 gpc1_1_5079(
      {stage059[140]},
      {stage059[233]}
   );
   gpc1_1 gpc1_1_5080(
      {stage059[141]},
      {stage059[234]}
   );
   gpc1_1 gpc1_1_5081(
      {stage059[142]},
      {stage059[235]}
   );
   gpc1_1 gpc1_1_5082(
      {stage059[143]},
      {stage059[236]}
   );
   gpc1_1 gpc1_1_5083(
      {stage059[144]},
      {stage059[237]}
   );
   gpc1_1 gpc1_1_5084(
      {stage059[145]},
      {stage059[238]}
   );
   gpc1_1 gpc1_1_5085(
      {stage059[146]},
      {stage059[239]}
   );
   gpc1_1 gpc1_1_5086(
      {stage059[147]},
      {stage059[240]}
   );
   gpc1_1 gpc1_1_5087(
      {stage059[148]},
      {stage059[241]}
   );
   gpc1_1 gpc1_1_5088(
      {stage059[149]},
      {stage059[242]}
   );
   gpc1_1 gpc1_1_5089(
      {stage059[150]},
      {stage059[243]}
   );
   gpc1_1 gpc1_1_5090(
      {stage059[151]},
      {stage059[244]}
   );
   gpc1_1 gpc1_1_5091(
      {stage059[152]},
      {stage059[245]}
   );
   gpc1_1 gpc1_1_5092(
      {stage059[153]},
      {stage059[246]}
   );
   gpc1_1 gpc1_1_5093(
      {stage059[154]},
      {stage059[247]}
   );
   gpc1_1 gpc1_1_5094(
      {stage059[155]},
      {stage059[248]}
   );
   gpc1_1 gpc1_1_5095(
      {stage059[156]},
      {stage059[249]}
   );
   gpc1_1 gpc1_1_5096(
      {stage059[157]},
      {stage059[250]}
   );
   gpc1_1 gpc1_1_5097(
      {stage059[158]},
      {stage059[251]}
   );
   gpc1_1 gpc1_1_5098(
      {stage059[159]},
      {stage059[252]}
   );
   gpc1_1 gpc1_1_5099(
      {stage059[160]},
      {stage059[253]}
   );
   gpc1_1 gpc1_1_5100(
      {stage059[161]},
      {stage059[254]}
   );
   gpc1_1 gpc1_1_5101(
      {stage059[162]},
      {stage059[255]}
   );
   gpc1_1 gpc1_1_5102(
      {stage059[163]},
      {stage059[256]}
   );
   gpc1_1 gpc1_1_5103(
      {stage059[164]},
      {stage059[257]}
   );
   gpc1_1 gpc1_1_5104(
      {stage059[165]},
      {stage059[258]}
   );
   gpc1_1 gpc1_1_5105(
      {stage059[166]},
      {stage059[259]}
   );
   gpc7_3 gpc7_3_5106(
      {stage059[167], stage059[168], stage059[169], stage059[170], stage059[171], stage059[172], stage059[173]},
      {stage061[197], stage060[199], stage059[260]}
   );
   gpc7_3 gpc7_3_5107(
      {stage059[174], stage059[175], stage059[176], stage059[177], stage059[178], stage059[179], stage059[180]},
      {stage061[198], stage060[200], stage059[261]}
   );
   gpc7_3 gpc7_3_5108(
      {stage059[181], stage059[182], stage059[183], stage059[184], stage059[185], stage059[186], stage059[187]},
      {stage061[199], stage060[201], stage059[262]}
   );
   gpc7_3 gpc7_3_5109(
      {stage059[188], stage059[189], stage059[190], stage059[191], stage059[192], stage059[193], stage059[194]},
      {stage061[200], stage060[202], stage059[263]}
   );
   gpc7_3 gpc7_3_5110(
      {stage059[195], stage059[196], stage059[197], stage059[198], stage059[199], stage059[200], stage059[201]},
      {stage061[201], stage060[203], stage059[264]}
   );
   gpc7_3 gpc7_3_5111(
      {stage059[202], stage059[203], stage059[204], stage059[205], stage059[206], stage059[207], stage059[208]},
      {stage061[202], stage060[204], stage059[265]}
   );
   gpc7_3 gpc7_3_5112(
      {stage059[209], stage059[210], stage059[211], stage059[212], stage059[213], stage059[214], stage059[215]},
      {stage061[203], stage060[205], stage059[266]}
   );
   gpc1_1 gpc1_1_5113(
      {stage060[176]},
      {stage060[206]}
   );
   gpc1_1 gpc1_1_5114(
      {stage060[177]},
      {stage060[207]}
   );
   gpc1_1 gpc1_1_5115(
      {stage060[178]},
      {stage060[208]}
   );
   gpc1_1 gpc1_1_5116(
      {stage060[179]},
      {stage060[209]}
   );
   gpc1_1 gpc1_1_5117(
      {stage060[180]},
      {stage060[210]}
   );
   gpc1_1 gpc1_1_5118(
      {stage060[181]},
      {stage060[211]}
   );
   gpc1_1 gpc1_1_5119(
      {stage060[182]},
      {stage060[212]}
   );
   gpc1_1 gpc1_1_5120(
      {stage060[183]},
      {stage060[213]}
   );
   gpc606_5 gpc606_5_5121(
      {stage060[184], stage060[185], stage060[186], stage060[187], stage060[188], stage060[189]},
      {stage062[128], stage062[129], stage062[130], stage062[131], stage062[132], stage062[133]},
      {stage064[211], stage063[175], stage062[197], stage061[204], stage060[214]}
   );
   gpc1_1 gpc1_1_5122(
      {stage061[128]},
      {stage061[205]}
   );
   gpc1_1 gpc1_1_5123(
      {stage061[129]},
      {stage061[206]}
   );
   gpc1_1 gpc1_1_5124(
      {stage061[130]},
      {stage061[207]}
   );
   gpc1_1 gpc1_1_5125(
      {stage061[131]},
      {stage061[208]}
   );
   gpc1_1 gpc1_1_5126(
      {stage061[132]},
      {stage061[209]}
   );
   gpc1_1 gpc1_1_5127(
      {stage061[133]},
      {stage061[210]}
   );
   gpc1_1 gpc1_1_5128(
      {stage061[134]},
      {stage061[211]}
   );
   gpc1_1 gpc1_1_5129(
      {stage061[135]},
      {stage061[212]}
   );
   gpc1_1 gpc1_1_5130(
      {stage061[136]},
      {stage061[213]}
   );
   gpc1_1 gpc1_1_5131(
      {stage061[137]},
      {stage061[214]}
   );
   gpc1_1 gpc1_1_5132(
      {stage061[138]},
      {stage061[215]}
   );
   gpc1_1 gpc1_1_5133(
      {stage061[139]},
      {stage061[216]}
   );
   gpc1_1 gpc1_1_5134(
      {stage061[140]},
      {stage061[217]}
   );
   gpc1_1 gpc1_1_5135(
      {stage061[141]},
      {stage061[218]}
   );
   gpc1_1 gpc1_1_5136(
      {stage061[142]},
      {stage061[219]}
   );
   gpc1_1 gpc1_1_5137(
      {stage061[143]},
      {stage061[220]}
   );
   gpc1_1 gpc1_1_5138(
      {stage061[144]},
      {stage061[221]}
   );
   gpc1_1 gpc1_1_5139(
      {stage061[145]},
      {stage061[222]}
   );
   gpc1_1 gpc1_1_5140(
      {stage061[146]},
      {stage061[223]}
   );
   gpc1_1 gpc1_1_5141(
      {stage061[147]},
      {stage061[224]}
   );
   gpc1_1 gpc1_1_5142(
      {stage061[148]},
      {stage061[225]}
   );
   gpc1_1 gpc1_1_5143(
      {stage061[149]},
      {stage061[226]}
   );
   gpc1_1 gpc1_1_5144(
      {stage061[150]},
      {stage061[227]}
   );
   gpc1_1 gpc1_1_5145(
      {stage061[151]},
      {stage061[228]}
   );
   gpc1_1 gpc1_1_5146(
      {stage061[152]},
      {stage061[229]}
   );
   gpc1_1 gpc1_1_5147(
      {stage061[153]},
      {stage061[230]}
   );
   gpc1_1 gpc1_1_5148(
      {stage061[154]},
      {stage061[231]}
   );
   gpc1_1 gpc1_1_5149(
      {stage061[155]},
      {stage061[232]}
   );
   gpc1_1 gpc1_1_5150(
      {stage061[156]},
      {stage061[233]}
   );
   gpc1_1 gpc1_1_5151(
      {stage061[157]},
      {stage061[234]}
   );
   gpc1_1 gpc1_1_5152(
      {stage061[158]},
      {stage061[235]}
   );
   gpc1_1 gpc1_1_5153(
      {stage061[159]},
      {stage061[236]}
   );
   gpc1_1 gpc1_1_5154(
      {stage061[160]},
      {stage061[237]}
   );
   gpc1_1 gpc1_1_5155(
      {stage061[161]},
      {stage061[238]}
   );
   gpc1_1 gpc1_1_5156(
      {stage061[162]},
      {stage061[239]}
   );
   gpc1_1 gpc1_1_5157(
      {stage061[163]},
      {stage061[240]}
   );
   gpc1_1 gpc1_1_5158(
      {stage061[164]},
      {stage061[241]}
   );
   gpc606_5 gpc606_5_5159(
      {stage061[165], stage061[166], stage061[167], stage061[168], stage061[169], stage061[170]},
      {stage063[128], stage063[129], stage063[130], stage063[131], stage063[132], stage063[133]},
      {stage065[199], stage064[212], stage063[176], stage062[198], stage061[242]}
   );
   gpc606_5 gpc606_5_5160(
      {stage061[171], stage061[172], stage061[173], stage061[174], stage061[175], stage061[176]},
      {stage063[134], stage063[135], stage063[136], stage063[137], stage063[138], stage063[139]},
      {stage065[200], stage064[213], stage063[177], stage062[199], stage061[243]}
   );
   gpc606_5 gpc606_5_5161(
      {stage061[177], stage061[178], stage061[179], stage061[180], stage061[181], stage061[182]},
      {stage063[140], stage063[141], stage063[142], stage063[143], stage063[144], stage063[145]},
      {stage065[201], stage064[214], stage063[178], stage062[200], stage061[244]}
   );
   gpc606_5 gpc606_5_5162(
      {stage061[183], stage061[184], stage061[185], stage061[186], stage061[187], stage061[188]},
      {stage063[146], stage063[147], stage063[148], stage063[149], stage063[150], stage063[151]},
      {stage065[202], stage064[215], stage063[179], stage062[201], stage061[245]}
   );
   gpc1_1 gpc1_1_5163(
      {stage062[134]},
      {stage062[202]}
   );
   gpc1_1 gpc1_1_5164(
      {stage062[135]},
      {stage062[203]}
   );
   gpc1_1 gpc1_1_5165(
      {stage062[136]},
      {stage062[204]}
   );
   gpc1_1 gpc1_1_5166(
      {stage062[137]},
      {stage062[205]}
   );
   gpc606_5 gpc606_5_5167(
      {stage062[138], stage062[139], stage062[140], stage062[141], stage062[142], stage062[143]},
      {stage064[128], stage064[129], stage064[130], stage064[131], stage064[132], stage064[133]},
      {stage066[211], stage065[203], stage064[216], stage063[180], stage062[206]}
   );
   gpc606_5 gpc606_5_5168(
      {stage062[144], stage062[145], stage062[146], stage062[147], stage062[148], stage062[149]},
      {stage064[134], stage064[135], stage064[136], stage064[137], stage064[138], stage064[139]},
      {stage066[212], stage065[204], stage064[217], stage063[181], stage062[207]}
   );
   gpc606_5 gpc606_5_5169(
      {stage062[150], stage062[151], stage062[152], stage062[153], stage062[154], stage062[155]},
      {stage064[140], stage064[141], stage064[142], stage064[143], stage064[144], stage064[145]},
      {stage066[213], stage065[205], stage064[218], stage063[182], stage062[208]}
   );
   gpc606_5 gpc606_5_5170(
      {stage062[156], stage062[157], stage062[158], stage062[159], stage062[160], stage062[161]},
      {stage064[146], stage064[147], stage064[148], stage064[149], stage064[150], stage064[151]},
      {stage066[214], stage065[206], stage064[219], stage063[183], stage062[209]}
   );
   gpc606_5 gpc606_5_5171(
      {stage062[162], stage062[163], stage062[164], stage062[165], stage062[166], stage062[167]},
      {stage064[152], stage064[153], stage064[154], stage064[155], stage064[156], stage064[157]},
      {stage066[215], stage065[207], stage064[220], stage063[184], stage062[210]}
   );
   gpc606_5 gpc606_5_5172(
      {stage062[168], stage062[169], stage062[170], stage062[171], stage062[172], stage062[173]},
      {stage064[158], stage064[159], stage064[160], stage064[161], stage064[162], stage064[163]},
      {stage066[216], stage065[208], stage064[221], stage063[185], stage062[211]}
   );
   gpc615_5 gpc615_5_5173(
      {stage062[174], stage062[175], stage062[176], stage062[177], stage062[178]},
      {stage063[152]},
      {stage064[164], stage064[165], stage064[166], stage064[167], stage064[168], stage064[169]},
      {stage066[217], stage065[209], stage064[222], stage063[186], stage062[212]}
   );
   gpc615_5 gpc615_5_5174(
      {stage062[179], stage062[180], stage062[181], stage062[182], stage062[183]},
      {stage063[153]},
      {stage064[170], stage064[171], stage064[172], stage064[173], stage064[174], stage064[175]},
      {stage066[218], stage065[210], stage064[223], stage063[187], stage062[213]}
   );
   gpc615_5 gpc615_5_5175(
      {stage062[184], stage062[185], stage062[186], stage062[187], stage062[188]},
      {stage063[154]},
      {stage064[176], stage064[177], stage064[178], stage064[179], stage064[180], stage064[181]},
      {stage066[219], stage065[211], stage064[224], stage063[188], stage062[214]}
   );
   gpc615_5 gpc615_5_5176(
      {stage063[155], stage063[156], stage063[157], stage063[158], stage063[159]},
      {stage064[182]},
      {stage065[128], stage065[129], stage065[130], stage065[131], stage065[132], stage065[133]},
      {stage067[213], stage066[220], stage065[212], stage064[225], stage063[189]}
   );
   gpc615_5 gpc615_5_5177(
      {stage063[160], stage063[161], stage063[162], stage063[163], stage063[164]},
      {stage064[183]},
      {stage065[134], stage065[135], stage065[136], stage065[137], stage065[138], stage065[139]},
      {stage067[214], stage066[221], stage065[213], stage064[226], stage063[190]}
   );
   gpc615_5 gpc615_5_5178(
      {stage063[165], stage063[166], stage063[167], stage063[168], stage063[169]},
      {stage064[184]},
      {stage065[140], stage065[141], stage065[142], stage065[143], stage065[144], stage065[145]},
      {stage067[215], stage066[222], stage065[214], stage064[227], stage063[191]}
   );
   gpc615_5 gpc615_5_5179(
      {stage063[170], stage063[171], stage063[172], stage063[173], stage063[174]},
      {stage064[185]},
      {stage065[146], stage065[147], stage065[148], stage065[149], stage065[150], stage065[151]},
      {stage067[216], stage066[223], stage065[215], stage064[228], stage063[192]}
   );
   gpc1_1 gpc1_1_5180(
      {stage064[186]},
      {stage064[229]}
   );
   gpc1_1 gpc1_1_5181(
      {stage064[187]},
      {stage064[230]}
   );
   gpc1_1 gpc1_1_5182(
      {stage064[188]},
      {stage064[231]}
   );
   gpc1_1 gpc1_1_5183(
      {stage064[189]},
      {stage064[232]}
   );
   gpc1_1 gpc1_1_5184(
      {stage064[190]},
      {stage064[233]}
   );
   gpc1_1 gpc1_1_5185(
      {stage064[191]},
      {stage064[234]}
   );
   gpc1_1 gpc1_1_5186(
      {stage064[192]},
      {stage064[235]}
   );
   gpc1_1 gpc1_1_5187(
      {stage064[193]},
      {stage064[236]}
   );
   gpc1_1 gpc1_1_5188(
      {stage064[194]},
      {stage064[237]}
   );
   gpc1_1 gpc1_1_5189(
      {stage064[195]},
      {stage064[238]}
   );
   gpc1_1 gpc1_1_5190(
      {stage064[196]},
      {stage064[239]}
   );
   gpc1_1 gpc1_1_5191(
      {stage064[197]},
      {stage064[240]}
   );
   gpc1_1 gpc1_1_5192(
      {stage064[198]},
      {stage064[241]}
   );
   gpc606_5 gpc606_5_5193(
      {stage064[199], stage064[200], stage064[201], stage064[202], stage064[203], stage064[204]},
      {stage066[128], stage066[129], stage066[130], stage066[131], stage066[132], stage066[133]},
      {stage068[210], stage067[217], stage066[224], stage065[216], stage064[242]}
   );
   gpc606_5 gpc606_5_5194(
      {stage064[205], stage064[206], stage064[207], stage064[208], stage064[209], stage064[210]},
      {stage066[134], stage066[135], stage066[136], stage066[137], stage066[138], stage066[139]},
      {stage068[211], stage067[218], stage066[225], stage065[217], stage064[243]}
   );
   gpc1_1 gpc1_1_5195(
      {stage065[152]},
      {stage065[218]}
   );
   gpc1_1 gpc1_1_5196(
      {stage065[153]},
      {stage065[219]}
   );
   gpc1_1 gpc1_1_5197(
      {stage065[154]},
      {stage065[220]}
   );
   gpc1_1 gpc1_1_5198(
      {stage065[155]},
      {stage065[221]}
   );
   gpc1_1 gpc1_1_5199(
      {stage065[156]},
      {stage065[222]}
   );
   gpc1_1 gpc1_1_5200(
      {stage065[157]},
      {stage065[223]}
   );
   gpc1_1 gpc1_1_5201(
      {stage065[158]},
      {stage065[224]}
   );
   gpc1_1 gpc1_1_5202(
      {stage065[159]},
      {stage065[225]}
   );
   gpc1_1 gpc1_1_5203(
      {stage065[160]},
      {stage065[226]}
   );
   gpc1_1 gpc1_1_5204(
      {stage065[161]},
      {stage065[227]}
   );
   gpc1_1 gpc1_1_5205(
      {stage065[162]},
      {stage065[228]}
   );
   gpc1_1 gpc1_1_5206(
      {stage065[163]},
      {stage065[229]}
   );
   gpc615_5 gpc615_5_5207(
      {stage065[164], stage065[165], stage065[166], stage065[167], stage065[168]},
      {stage066[140]},
      {stage067[128], stage067[129], stage067[130], stage067[131], stage067[132], stage067[133]},
      {stage069[183], stage068[212], stage067[219], stage066[226], stage065[230]}
   );
   gpc615_5 gpc615_5_5208(
      {stage065[169], stage065[170], stage065[171], stage065[172], stage065[173]},
      {stage066[141]},
      {stage067[134], stage067[135], stage067[136], stage067[137], stage067[138], stage067[139]},
      {stage069[184], stage068[213], stage067[220], stage066[227], stage065[231]}
   );
   gpc615_5 gpc615_5_5209(
      {stage065[174], stage065[175], stage065[176], stage065[177], stage065[178]},
      {stage066[142]},
      {stage067[140], stage067[141], stage067[142], stage067[143], stage067[144], stage067[145]},
      {stage069[185], stage068[214], stage067[221], stage066[228], stage065[232]}
   );
   gpc615_5 gpc615_5_5210(
      {stage065[179], stage065[180], stage065[181], stage065[182], stage065[183]},
      {stage066[143]},
      {stage067[146], stage067[147], stage067[148], stage067[149], stage067[150], stage067[151]},
      {stage069[186], stage068[215], stage067[222], stage066[229], stage065[233]}
   );
   gpc615_5 gpc615_5_5211(
      {stage065[184], stage065[185], stage065[186], stage065[187], stage065[188]},
      {stage066[144]},
      {stage067[152], stage067[153], stage067[154], stage067[155], stage067[156], stage067[157]},
      {stage069[187], stage068[216], stage067[223], stage066[230], stage065[234]}
   );
   gpc615_5 gpc615_5_5212(
      {stage065[189], stage065[190], stage065[191], stage065[192], stage065[193]},
      {stage066[145]},
      {stage067[158], stage067[159], stage067[160], stage067[161], stage067[162], stage067[163]},
      {stage069[188], stage068[217], stage067[224], stage066[231], stage065[235]}
   );
   gpc615_5 gpc615_5_5213(
      {stage065[194], stage065[195], stage065[196], stage065[197], stage065[198]},
      {stage066[146]},
      {stage067[164], stage067[165], stage067[166], stage067[167], stage067[168], stage067[169]},
      {stage069[189], stage068[218], stage067[225], stage066[232], stage065[236]}
   );
   gpc615_5 gpc615_5_5214(
      {stage066[147], stage066[148], stage066[149], stage066[150], stage066[151]},
      {stage067[170]},
      {stage068[128], stage068[129], stage068[130], stage068[131], stage068[132], stage068[133]},
      {stage070[189], stage069[190], stage068[219], stage067[226], stage066[233]}
   );
   gpc615_5 gpc615_5_5215(
      {stage066[152], stage066[153], stage066[154], stage066[155], stage066[156]},
      {stage067[171]},
      {stage068[134], stage068[135], stage068[136], stage068[137], stage068[138], stage068[139]},
      {stage070[190], stage069[191], stage068[220], stage067[227], stage066[234]}
   );
   gpc615_5 gpc615_5_5216(
      {stage066[157], stage066[158], stage066[159], stage066[160], stage066[161]},
      {stage067[172]},
      {stage068[140], stage068[141], stage068[142], stage068[143], stage068[144], stage068[145]},
      {stage070[191], stage069[192], stage068[221], stage067[228], stage066[235]}
   );
   gpc615_5 gpc615_5_5217(
      {stage066[162], stage066[163], stage066[164], stage066[165], stage066[166]},
      {stage067[173]},
      {stage068[146], stage068[147], stage068[148], stage068[149], stage068[150], stage068[151]},
      {stage070[192], stage069[193], stage068[222], stage067[229], stage066[236]}
   );
   gpc615_5 gpc615_5_5218(
      {stage066[167], stage066[168], stage066[169], stage066[170], stage066[171]},
      {stage067[174]},
      {stage068[152], stage068[153], stage068[154], stage068[155], stage068[156], stage068[157]},
      {stage070[193], stage069[194], stage068[223], stage067[230], stage066[237]}
   );
   gpc615_5 gpc615_5_5219(
      {stage066[172], stage066[173], stage066[174], stage066[175], stage066[176]},
      {stage067[175]},
      {stage068[158], stage068[159], stage068[160], stage068[161], stage068[162], stage068[163]},
      {stage070[194], stage069[195], stage068[224], stage067[231], stage066[238]}
   );
   gpc615_5 gpc615_5_5220(
      {stage066[177], stage066[178], stage066[179], stage066[180], stage066[181]},
      {stage067[176]},
      {stage068[164], stage068[165], stage068[166], stage068[167], stage068[168], stage068[169]},
      {stage070[195], stage069[196], stage068[225], stage067[232], stage066[239]}
   );
   gpc615_5 gpc615_5_5221(
      {stage066[182], stage066[183], stage066[184], stage066[185], stage066[186]},
      {stage067[177]},
      {stage068[170], stage068[171], stage068[172], stage068[173], stage068[174], stage068[175]},
      {stage070[196], stage069[197], stage068[226], stage067[233], stage066[240]}
   );
   gpc615_5 gpc615_5_5222(
      {stage066[187], stage066[188], stage066[189], stage066[190], stage066[191]},
      {stage067[178]},
      {stage068[176], stage068[177], stage068[178], stage068[179], stage068[180], stage068[181]},
      {stage070[197], stage069[198], stage068[227], stage067[234], stage066[241]}
   );
   gpc615_5 gpc615_5_5223(
      {stage066[192], stage066[193], stage066[194], stage066[195], stage066[196]},
      {stage067[179]},
      {stage068[182], stage068[183], stage068[184], stage068[185], stage068[186], stage068[187]},
      {stage070[198], stage069[199], stage068[228], stage067[235], stage066[242]}
   );
   gpc615_5 gpc615_5_5224(
      {stage066[197], stage066[198], stage066[199], stage066[200], stage066[201]},
      {stage067[180]},
      {stage068[188], stage068[189], stage068[190], stage068[191], stage068[192], stage068[193]},
      {stage070[199], stage069[200], stage068[229], stage067[236], stage066[243]}
   );
   gpc615_5 gpc615_5_5225(
      {stage066[202], stage066[203], stage066[204], stage066[205], stage066[206]},
      {stage067[181]},
      {stage068[194], stage068[195], stage068[196], stage068[197], stage068[198], stage068[199]},
      {stage070[200], stage069[201], stage068[230], stage067[237], stage066[244]}
   );
   gpc615_5 gpc615_5_5226(
      {stage066[207], stage066[208], stage066[209], stage066[210], 1'h0},
      {stage067[182]},
      {stage068[200], stage068[201], stage068[202], stage068[203], stage068[204], stage068[205]},
      {stage070[201], stage069[202], stage068[231], stage067[238], stage066[245]}
   );
   gpc606_5 gpc606_5_5227(
      {stage067[183], stage067[184], stage067[185], stage067[186], stage067[187], stage067[188]},
      {stage069[128], stage069[129], stage069[130], stage069[131], stage069[132], stage069[133]},
      {stage071[188], stage070[202], stage069[203], stage068[232], stage067[239]}
   );
   gpc606_5 gpc606_5_5228(
      {stage067[189], stage067[190], stage067[191], stage067[192], stage067[193], stage067[194]},
      {stage069[134], stage069[135], stage069[136], stage069[137], stage069[138], stage069[139]},
      {stage071[189], stage070[203], stage069[204], stage068[233], stage067[240]}
   );
   gpc606_5 gpc606_5_5229(
      {stage067[195], stage067[196], stage067[197], stage067[198], stage067[199], stage067[200]},
      {stage069[140], stage069[141], stage069[142], stage069[143], stage069[144], stage069[145]},
      {stage071[190], stage070[204], stage069[205], stage068[234], stage067[241]}
   );
   gpc606_5 gpc606_5_5230(
      {stage067[201], stage067[202], stage067[203], stage067[204], stage067[205], stage067[206]},
      {stage069[146], stage069[147], stage069[148], stage069[149], stage069[150], stage069[151]},
      {stage071[191], stage070[205], stage069[206], stage068[235], stage067[242]}
   );
   gpc606_5 gpc606_5_5231(
      {stage067[207], stage067[208], stage067[209], stage067[210], stage067[211], stage067[212]},
      {stage069[152], stage069[153], stage069[154], stage069[155], stage069[156], stage069[157]},
      {stage071[192], stage070[206], stage069[207], stage068[236], stage067[243]}
   );
   gpc1_1 gpc1_1_5232(
      {stage068[206]},
      {stage068[237]}
   );
   gpc1_1 gpc1_1_5233(
      {stage068[207]},
      {stage068[238]}
   );
   gpc1_1 gpc1_1_5234(
      {stage068[208]},
      {stage068[239]}
   );
   gpc1_1 gpc1_1_5235(
      {stage068[209]},
      {stage068[240]}
   );
   gpc1_1 gpc1_1_5236(
      {stage069[158]},
      {stage069[208]}
   );
   gpc1_1 gpc1_1_5237(
      {stage069[159]},
      {stage069[209]}
   );
   gpc1_1 gpc1_1_5238(
      {stage069[160]},
      {stage069[210]}
   );
   gpc1_1 gpc1_1_5239(
      {stage069[161]},
      {stage069[211]}
   );
   gpc1_1 gpc1_1_5240(
      {stage069[162]},
      {stage069[212]}
   );
   gpc1_1 gpc1_1_5241(
      {stage069[163]},
      {stage069[213]}
   );
   gpc1_1 gpc1_1_5242(
      {stage069[164]},
      {stage069[214]}
   );
   gpc1_1 gpc1_1_5243(
      {stage069[165]},
      {stage069[215]}
   );
   gpc1_1 gpc1_1_5244(
      {stage069[166]},
      {stage069[216]}
   );
   gpc1_1 gpc1_1_5245(
      {stage069[167]},
      {stage069[217]}
   );
   gpc1_1 gpc1_1_5246(
      {stage069[168]},
      {stage069[218]}
   );
   gpc1_1 gpc1_1_5247(
      {stage069[169]},
      {stage069[219]}
   );
   gpc1_1 gpc1_1_5248(
      {stage069[170]},
      {stage069[220]}
   );
   gpc1_1 gpc1_1_5249(
      {stage069[171]},
      {stage069[221]}
   );
   gpc1_1 gpc1_1_5250(
      {stage069[172]},
      {stage069[222]}
   );
   gpc1_1 gpc1_1_5251(
      {stage069[173]},
      {stage069[223]}
   );
   gpc1_1 gpc1_1_5252(
      {stage069[174]},
      {stage069[224]}
   );
   gpc1_1 gpc1_1_5253(
      {stage069[175]},
      {stage069[225]}
   );
   gpc1_1 gpc1_1_5254(
      {stage069[176]},
      {stage069[226]}
   );
   gpc1_1 gpc1_1_5255(
      {stage069[177]},
      {stage069[227]}
   );
   gpc1_1 gpc1_1_5256(
      {stage069[178]},
      {stage069[228]}
   );
   gpc1_1 gpc1_1_5257(
      {stage069[179]},
      {stage069[229]}
   );
   gpc1_1 gpc1_1_5258(
      {stage069[180]},
      {stage069[230]}
   );
   gpc1_1 gpc1_1_5259(
      {stage069[181]},
      {stage069[231]}
   );
   gpc1_1 gpc1_1_5260(
      {stage069[182]},
      {stage069[232]}
   );
   gpc1_1 gpc1_1_5261(
      {stage070[128]},
      {stage070[207]}
   );
   gpc1_1 gpc1_1_5262(
      {stage070[129]},
      {stage070[208]}
   );
   gpc1_1 gpc1_1_5263(
      {stage070[130]},
      {stage070[209]}
   );
   gpc1_1 gpc1_1_5264(
      {stage070[131]},
      {stage070[210]}
   );
   gpc1_1 gpc1_1_5265(
      {stage070[132]},
      {stage070[211]}
   );
   gpc1_1 gpc1_1_5266(
      {stage070[133]},
      {stage070[212]}
   );
   gpc1_1 gpc1_1_5267(
      {stage070[134]},
      {stage070[213]}
   );
   gpc1_1 gpc1_1_5268(
      {stage070[135]},
      {stage070[214]}
   );
   gpc1_1 gpc1_1_5269(
      {stage070[136]},
      {stage070[215]}
   );
   gpc1_1 gpc1_1_5270(
      {stage070[137]},
      {stage070[216]}
   );
   gpc1_1 gpc1_1_5271(
      {stage070[138]},
      {stage070[217]}
   );
   gpc1_1 gpc1_1_5272(
      {stage070[139]},
      {stage070[218]}
   );
   gpc1_1 gpc1_1_5273(
      {stage070[140]},
      {stage070[219]}
   );
   gpc1_1 gpc1_1_5274(
      {stage070[141]},
      {stage070[220]}
   );
   gpc1_1 gpc1_1_5275(
      {stage070[142]},
      {stage070[221]}
   );
   gpc1_1 gpc1_1_5276(
      {stage070[143]},
      {stage070[222]}
   );
   gpc1_1 gpc1_1_5277(
      {stage070[144]},
      {stage070[223]}
   );
   gpc1_1 gpc1_1_5278(
      {stage070[145]},
      {stage070[224]}
   );
   gpc1_1 gpc1_1_5279(
      {stage070[146]},
      {stage070[225]}
   );
   gpc606_5 gpc606_5_5280(
      {stage070[147], stage070[148], stage070[149], stage070[150], stage070[151], stage070[152]},
      {stage072[128], stage072[129], stage072[130], stage072[131], stage072[132], stage072[133]},
      {stage074[189], stage073[193], stage072[222], stage071[193], stage070[226]}
   );
   gpc606_5 gpc606_5_5281(
      {stage070[153], stage070[154], stage070[155], stage070[156], stage070[157], stage070[158]},
      {stage072[134], stage072[135], stage072[136], stage072[137], stage072[138], stage072[139]},
      {stage074[190], stage073[194], stage072[223], stage071[194], stage070[227]}
   );
   gpc615_5 gpc615_5_5282(
      {stage070[159], stage070[160], stage070[161], stage070[162], stage070[163]},
      {stage071[128]},
      {stage072[140], stage072[141], stage072[142], stage072[143], stage072[144], stage072[145]},
      {stage074[191], stage073[195], stage072[224], stage071[195], stage070[228]}
   );
   gpc615_5 gpc615_5_5283(
      {stage070[164], stage070[165], stage070[166], stage070[167], stage070[168]},
      {stage071[129]},
      {stage072[146], stage072[147], stage072[148], stage072[149], stage072[150], stage072[151]},
      {stage074[192], stage073[196], stage072[225], stage071[196], stage070[229]}
   );
   gpc615_5 gpc615_5_5284(
      {stage070[169], stage070[170], stage070[171], stage070[172], stage070[173]},
      {stage071[130]},
      {stage072[152], stage072[153], stage072[154], stage072[155], stage072[156], stage072[157]},
      {stage074[193], stage073[197], stage072[226], stage071[197], stage070[230]}
   );
   gpc615_5 gpc615_5_5285(
      {stage070[174], stage070[175], stage070[176], stage070[177], stage070[178]},
      {stage071[131]},
      {stage072[158], stage072[159], stage072[160], stage072[161], stage072[162], stage072[163]},
      {stage074[194], stage073[198], stage072[227], stage071[198], stage070[231]}
   );
   gpc615_5 gpc615_5_5286(
      {stage070[179], stage070[180], stage070[181], stage070[182], stage070[183]},
      {stage071[132]},
      {stage072[164], stage072[165], stage072[166], stage072[167], stage072[168], stage072[169]},
      {stage074[195], stage073[199], stage072[228], stage071[199], stage070[232]}
   );
   gpc615_5 gpc615_5_5287(
      {stage070[184], stage070[185], stage070[186], stage070[187], stage070[188]},
      {stage071[133]},
      {stage072[170], stage072[171], stage072[172], stage072[173], stage072[174], stage072[175]},
      {stage074[196], stage073[200], stage072[229], stage071[200], stage070[233]}
   );
   gpc1_1 gpc1_1_5288(
      {stage071[134]},
      {stage071[201]}
   );
   gpc1_1 gpc1_1_5289(
      {stage071[135]},
      {stage071[202]}
   );
   gpc1_1 gpc1_1_5290(
      {stage071[136]},
      {stage071[203]}
   );
   gpc1_1 gpc1_1_5291(
      {stage071[137]},
      {stage071[204]}
   );
   gpc1_1 gpc1_1_5292(
      {stage071[138]},
      {stage071[205]}
   );
   gpc1_1 gpc1_1_5293(
      {stage071[139]},
      {stage071[206]}
   );
   gpc1_1 gpc1_1_5294(
      {stage071[140]},
      {stage071[207]}
   );
   gpc1_1 gpc1_1_5295(
      {stage071[141]},
      {stage071[208]}
   );
   gpc1_1 gpc1_1_5296(
      {stage071[142]},
      {stage071[209]}
   );
   gpc1_1 gpc1_1_5297(
      {stage071[143]},
      {stage071[210]}
   );
   gpc1_1 gpc1_1_5298(
      {stage071[144]},
      {stage071[211]}
   );
   gpc1_1 gpc1_1_5299(
      {stage071[145]},
      {stage071[212]}
   );
   gpc1_1 gpc1_1_5300(
      {stage071[146]},
      {stage071[213]}
   );
   gpc1_1 gpc1_1_5301(
      {stage071[147]},
      {stage071[214]}
   );
   gpc1_1 gpc1_1_5302(
      {stage071[148]},
      {stage071[215]}
   );
   gpc1_1 gpc1_1_5303(
      {stage071[149]},
      {stage071[216]}
   );
   gpc1_1 gpc1_1_5304(
      {stage071[150]},
      {stage071[217]}
   );
   gpc1_1 gpc1_1_5305(
      {stage071[151]},
      {stage071[218]}
   );
   gpc1_1 gpc1_1_5306(
      {stage071[152]},
      {stage071[219]}
   );
   gpc1_1 gpc1_1_5307(
      {stage071[153]},
      {stage071[220]}
   );
   gpc1_1 gpc1_1_5308(
      {stage071[154]},
      {stage071[221]}
   );
   gpc1_1 gpc1_1_5309(
      {stage071[155]},
      {stage071[222]}
   );
   gpc1_1 gpc1_1_5310(
      {stage071[156]},
      {stage071[223]}
   );
   gpc1_1 gpc1_1_5311(
      {stage071[157]},
      {stage071[224]}
   );
   gpc1_1 gpc1_1_5312(
      {stage071[158]},
      {stage071[225]}
   );
   gpc1_1 gpc1_1_5313(
      {stage071[159]},
      {stage071[226]}
   );
   gpc1_1 gpc1_1_5314(
      {stage071[160]},
      {stage071[227]}
   );
   gpc623_5 gpc623_5_5315(
      {stage071[161], stage071[162], stage071[163]},
      {stage072[176], stage072[177]},
      {stage073[128], stage073[129], stage073[130], stage073[131], stage073[132], stage073[133]},
      {stage075[169], stage074[197], stage073[201], stage072[230], stage071[228]}
   );
   gpc623_5 gpc623_5_5316(
      {stage071[164], stage071[165], stage071[166]},
      {stage072[178], stage072[179]},
      {stage073[134], stage073[135], stage073[136], stage073[137], stage073[138], stage073[139]},
      {stage075[170], stage074[198], stage073[202], stage072[231], stage071[229]}
   );
   gpc623_5 gpc623_5_5317(
      {stage071[167], stage071[168], stage071[169]},
      {stage072[180], stage072[181]},
      {stage073[140], stage073[141], stage073[142], stage073[143], stage073[144], stage073[145]},
      {stage075[171], stage074[199], stage073[203], stage072[232], stage071[230]}
   );
   gpc623_5 gpc623_5_5318(
      {stage071[170], stage071[171], stage071[172]},
      {stage072[182], stage072[183]},
      {stage073[146], stage073[147], stage073[148], stage073[149], stage073[150], stage073[151]},
      {stage075[172], stage074[200], stage073[204], stage072[233], stage071[231]}
   );
   gpc623_5 gpc623_5_5319(
      {stage071[173], stage071[174], stage071[175]},
      {stage072[184], stage072[185]},
      {stage073[152], stage073[153], stage073[154], stage073[155], stage073[156], stage073[157]},
      {stage075[173], stage074[201], stage073[205], stage072[234], stage071[232]}
   );
   gpc623_5 gpc623_5_5320(
      {stage071[176], stage071[177], stage071[178]},
      {stage072[186], stage072[187]},
      {stage073[158], stage073[159], stage073[160], stage073[161], stage073[162], stage073[163]},
      {stage075[174], stage074[202], stage073[206], stage072[235], stage071[233]}
   );
   gpc623_5 gpc623_5_5321(
      {stage071[179], stage071[180], stage071[181]},
      {stage072[188], stage072[189]},
      {stage073[164], stage073[165], stage073[166], stage073[167], stage073[168], stage073[169]},
      {stage075[175], stage074[203], stage073[207], stage072[236], stage071[234]}
   );
   gpc623_5 gpc623_5_5322(
      {stage071[182], stage071[183], stage071[184]},
      {stage072[190], stage072[191]},
      {stage073[170], stage073[171], stage073[172], stage073[173], stage073[174], stage073[175]},
      {stage075[176], stage074[204], stage073[208], stage072[237], stage071[235]}
   );
   gpc623_5 gpc623_5_5323(
      {stage071[185], stage071[186], stage071[187]},
      {stage072[192], stage072[193]},
      {stage073[176], stage073[177], stage073[178], stage073[179], stage073[180], stage073[181]},
      {stage075[177], stage074[205], stage073[209], stage072[238], stage071[236]}
   );
   gpc1_1 gpc1_1_5324(
      {stage072[194]},
      {stage072[239]}
   );
   gpc1_1 gpc1_1_5325(
      {stage072[195]},
      {stage072[240]}
   );
   gpc1_1 gpc1_1_5326(
      {stage072[196]},
      {stage072[241]}
   );
   gpc1_1 gpc1_1_5327(
      {stage072[197]},
      {stage072[242]}
   );
   gpc1_1 gpc1_1_5328(
      {stage072[198]},
      {stage072[243]}
   );
   gpc1_1 gpc1_1_5329(
      {stage072[199]},
      {stage072[244]}
   );
   gpc1_1 gpc1_1_5330(
      {stage072[200]},
      {stage072[245]}
   );
   gpc1_1 gpc1_1_5331(
      {stage072[201]},
      {stage072[246]}
   );
   gpc1_1 gpc1_1_5332(
      {stage072[202]},
      {stage072[247]}
   );
   gpc1_1 gpc1_1_5333(
      {stage072[203]},
      {stage072[248]}
   );
   gpc1_1 gpc1_1_5334(
      {stage072[204]},
      {stage072[249]}
   );
   gpc1_1 gpc1_1_5335(
      {stage072[205]},
      {stage072[250]}
   );
   gpc1_1 gpc1_1_5336(
      {stage072[206]},
      {stage072[251]}
   );
   gpc1_1 gpc1_1_5337(
      {stage072[207]},
      {stage072[252]}
   );
   gpc1_1 gpc1_1_5338(
      {stage072[208]},
      {stage072[253]}
   );
   gpc1_1 gpc1_1_5339(
      {stage072[209]},
      {stage072[254]}
   );
   gpc1_1 gpc1_1_5340(
      {stage072[210]},
      {stage072[255]}
   );
   gpc1_1 gpc1_1_5341(
      {stage072[211]},
      {stage072[256]}
   );
   gpc1_1 gpc1_1_5342(
      {stage072[212]},
      {stage072[257]}
   );
   gpc1_1 gpc1_1_5343(
      {stage072[213]},
      {stage072[258]}
   );
   gpc1_1 gpc1_1_5344(
      {stage072[214]},
      {stage072[259]}
   );
   gpc1_1 gpc1_1_5345(
      {stage072[215]},
      {stage072[260]}
   );
   gpc1_1 gpc1_1_5346(
      {stage072[216]},
      {stage072[261]}
   );
   gpc1_1 gpc1_1_5347(
      {stage072[217]},
      {stage072[262]}
   );
   gpc1_1 gpc1_1_5348(
      {stage072[218]},
      {stage072[263]}
   );
   gpc1_1 gpc1_1_5349(
      {stage072[219]},
      {stage072[264]}
   );
   gpc1_1 gpc1_1_5350(
      {stage072[220]},
      {stage072[265]}
   );
   gpc1_1 gpc1_1_5351(
      {stage072[221]},
      {stage072[266]}
   );
   gpc1_1 gpc1_1_5352(
      {stage073[182]},
      {stage073[210]}
   );
   gpc1_1 gpc1_1_5353(
      {stage073[183]},
      {stage073[211]}
   );
   gpc1_1 gpc1_1_5354(
      {stage073[184]},
      {stage073[212]}
   );
   gpc1_1 gpc1_1_5355(
      {stage073[185]},
      {stage073[213]}
   );
   gpc1_1 gpc1_1_5356(
      {stage073[186]},
      {stage073[214]}
   );
   gpc1_1 gpc1_1_5357(
      {stage073[187]},
      {stage073[215]}
   );
   gpc615_5 gpc615_5_5358(
      {stage073[188], stage073[189], stage073[190], stage073[191], stage073[192]},
      {stage074[128]},
      {stage075[128], stage075[129], stage075[130], stage075[131], stage075[132], stage075[133]},
      {stage077[203], stage076[182], stage075[178], stage074[206], stage073[216]}
   );
   gpc1_1 gpc1_1_5359(
      {stage074[129]},
      {stage074[207]}
   );
   gpc1_1 gpc1_1_5360(
      {stage074[130]},
      {stage074[208]}
   );
   gpc1_1 gpc1_1_5361(
      {stage074[131]},
      {stage074[209]}
   );
   gpc1_1 gpc1_1_5362(
      {stage074[132]},
      {stage074[210]}
   );
   gpc1_1 gpc1_1_5363(
      {stage074[133]},
      {stage074[211]}
   );
   gpc1_1 gpc1_1_5364(
      {stage074[134]},
      {stage074[212]}
   );
   gpc1_1 gpc1_1_5365(
      {stage074[135]},
      {stage074[213]}
   );
   gpc1_1 gpc1_1_5366(
      {stage074[136]},
      {stage074[214]}
   );
   gpc1_1 gpc1_1_5367(
      {stage074[137]},
      {stage074[215]}
   );
   gpc1_1 gpc1_1_5368(
      {stage074[138]},
      {stage074[216]}
   );
   gpc1_1 gpc1_1_5369(
      {stage074[139]},
      {stage074[217]}
   );
   gpc606_5 gpc606_5_5370(
      {stage074[140], stage074[141], stage074[142], stage074[143], stage074[144], stage074[145]},
      {stage076[128], stage076[129], stage076[130], stage076[131], stage076[132], stage076[133]},
      {stage078[174], stage077[204], stage076[183], stage075[179], stage074[218]}
   );
   gpc606_5 gpc606_5_5371(
      {stage074[146], stage074[147], stage074[148], stage074[149], stage074[150], stage074[151]},
      {stage076[134], stage076[135], stage076[136], stage076[137], stage076[138], stage076[139]},
      {stage078[175], stage077[205], stage076[184], stage075[180], stage074[219]}
   );
   gpc606_5 gpc606_5_5372(
      {stage074[152], stage074[153], stage074[154], stage074[155], stage074[156], stage074[157]},
      {stage076[140], stage076[141], stage076[142], stage076[143], stage076[144], stage076[145]},
      {stage078[176], stage077[206], stage076[185], stage075[181], stage074[220]}
   );
   gpc606_5 gpc606_5_5373(
      {stage074[158], stage074[159], stage074[160], stage074[161], stage074[162], stage074[163]},
      {stage076[146], stage076[147], stage076[148], stage076[149], stage076[150], stage076[151]},
      {stage078[177], stage077[207], stage076[186], stage075[182], stage074[221]}
   );
   gpc615_5 gpc615_5_5374(
      {stage074[164], stage074[165], stage074[166], stage074[167], stage074[168]},
      {stage075[134]},
      {stage076[152], stage076[153], stage076[154], stage076[155], stage076[156], stage076[157]},
      {stage078[178], stage077[208], stage076[187], stage075[183], stage074[222]}
   );
   gpc615_5 gpc615_5_5375(
      {stage074[169], stage074[170], stage074[171], stage074[172], stage074[173]},
      {stage075[135]},
      {stage076[158], stage076[159], stage076[160], stage076[161], stage076[162], stage076[163]},
      {stage078[179], stage077[209], stage076[188], stage075[184], stage074[223]}
   );
   gpc615_5 gpc615_5_5376(
      {stage074[174], stage074[175], stage074[176], stage074[177], stage074[178]},
      {stage075[136]},
      {stage076[164], stage076[165], stage076[166], stage076[167], stage076[168], stage076[169]},
      {stage078[180], stage077[210], stage076[189], stage075[185], stage074[224]}
   );
   gpc615_5 gpc615_5_5377(
      {stage074[179], stage074[180], stage074[181], stage074[182], stage074[183]},
      {stage075[137]},
      {stage076[170], stage076[171], stage076[172], stage076[173], stage076[174], stage076[175]},
      {stage078[181], stage077[211], stage076[190], stage075[186], stage074[225]}
   );
   gpc615_5 gpc615_5_5378(
      {stage074[184], stage074[185], stage074[186], stage074[187], stage074[188]},
      {stage075[138]},
      {stage076[176], stage076[177], stage076[178], stage076[179], stage076[180], stage076[181]},
      {stage078[182], stage077[212], stage076[191], stage075[187], stage074[226]}
   );
   gpc606_5 gpc606_5_5379(
      {stage075[139], stage075[140], stage075[141], stage075[142], stage075[143], stage075[144]},
      {stage077[128], stage077[129], stage077[130], stage077[131], stage077[132], stage077[133]},
      {stage079[187], stage078[183], stage077[213], stage076[192], stage075[188]}
   );
   gpc606_5 gpc606_5_5380(
      {stage075[145], stage075[146], stage075[147], stage075[148], stage075[149], stage075[150]},
      {stage077[134], stage077[135], stage077[136], stage077[137], stage077[138], stage077[139]},
      {stage079[188], stage078[184], stage077[214], stage076[193], stage075[189]}
   );
   gpc606_5 gpc606_5_5381(
      {stage075[151], stage075[152], stage075[153], stage075[154], stage075[155], stage075[156]},
      {stage077[140], stage077[141], stage077[142], stage077[143], stage077[144], stage077[145]},
      {stage079[189], stage078[185], stage077[215], stage076[194], stage075[190]}
   );
   gpc606_5 gpc606_5_5382(
      {stage075[157], stage075[158], stage075[159], stage075[160], stage075[161], stage075[162]},
      {stage077[146], stage077[147], stage077[148], stage077[149], stage077[150], stage077[151]},
      {stage079[190], stage078[186], stage077[216], stage076[195], stage075[191]}
   );
   gpc606_5 gpc606_5_5383(
      {stage075[163], stage075[164], stage075[165], stage075[166], stage075[167], stage075[168]},
      {stage077[152], stage077[153], stage077[154], stage077[155], stage077[156], stage077[157]},
      {stage079[191], stage078[187], stage077[217], stage076[196], stage075[192]}
   );
   gpc1_1 gpc1_1_5384(
      {stage077[158]},
      {stage077[218]}
   );
   gpc1_1 gpc1_1_5385(
      {stage077[159]},
      {stage077[219]}
   );
   gpc1_1 gpc1_1_5386(
      {stage077[160]},
      {stage077[220]}
   );
   gpc1_1 gpc1_1_5387(
      {stage077[161]},
      {stage077[221]}
   );
   gpc1_1 gpc1_1_5388(
      {stage077[162]},
      {stage077[222]}
   );
   gpc606_5 gpc606_5_5389(
      {stage077[163], stage077[164], stage077[165], stage077[166], stage077[167], stage077[168]},
      {stage079[128], stage079[129], stage079[130], stage079[131], stage079[132], stage079[133]},
      {stage081[175], stage080[203], stage079[192], stage078[188], stage077[223]}
   );
   gpc606_5 gpc606_5_5390(
      {stage077[169], stage077[170], stage077[171], stage077[172], stage077[173], stage077[174]},
      {stage079[134], stage079[135], stage079[136], stage079[137], stage079[138], stage079[139]},
      {stage081[176], stage080[204], stage079[193], stage078[189], stage077[224]}
   );
   gpc606_5 gpc606_5_5391(
      {stage077[175], stage077[176], stage077[177], stage077[178], stage077[179], stage077[180]},
      {stage079[140], stage079[141], stage079[142], stage079[143], stage079[144], stage079[145]},
      {stage081[177], stage080[205], stage079[194], stage078[190], stage077[225]}
   );
   gpc606_5 gpc606_5_5392(
      {stage077[181], stage077[182], stage077[183], stage077[184], stage077[185], stage077[186]},
      {stage079[146], stage079[147], stage079[148], stage079[149], stage079[150], stage079[151]},
      {stage081[178], stage080[206], stage079[195], stage078[191], stage077[226]}
   );
   gpc606_5 gpc606_5_5393(
      {stage077[187], stage077[188], stage077[189], stage077[190], stage077[191], stage077[192]},
      {stage079[152], stage079[153], stage079[154], stage079[155], stage079[156], stage079[157]},
      {stage081[179], stage080[207], stage079[196], stage078[192], stage077[227]}
   );
   gpc615_5 gpc615_5_5394(
      {stage077[193], stage077[194], stage077[195], stage077[196], stage077[197]},
      {stage078[128]},
      {stage079[158], stage079[159], stage079[160], stage079[161], stage079[162], stage079[163]},
      {stage081[180], stage080[208], stage079[197], stage078[193], stage077[228]}
   );
   gpc615_5 gpc615_5_5395(
      {stage077[198], stage077[199], stage077[200], stage077[201], stage077[202]},
      {stage078[129]},
      {stage079[164], stage079[165], stage079[166], stage079[167], stage079[168], stage079[169]},
      {stage081[181], stage080[209], stage079[198], stage078[194], stage077[229]}
   );
   gpc1_1 gpc1_1_5396(
      {stage078[130]},
      {stage078[195]}
   );
   gpc1_1 gpc1_1_5397(
      {stage078[131]},
      {stage078[196]}
   );
   gpc1_1 gpc1_1_5398(
      {stage078[132]},
      {stage078[197]}
   );
   gpc1_1 gpc1_1_5399(
      {stage078[133]},
      {stage078[198]}
   );
   gpc615_5 gpc615_5_5400(
      {stage078[134], stage078[135], stage078[136], stage078[137], stage078[138]},
      {stage079[170]},
      {stage080[128], stage080[129], stage080[130], stage080[131], stage080[132], stage080[133]},
      {stage082[215], stage081[182], stage080[210], stage079[199], stage078[199]}
   );
   gpc615_5 gpc615_5_5401(
      {stage078[139], stage078[140], stage078[141], stage078[142], stage078[143]},
      {stage079[171]},
      {stage080[134], stage080[135], stage080[136], stage080[137], stage080[138], stage080[139]},
      {stage082[216], stage081[183], stage080[211], stage079[200], stage078[200]}
   );
   gpc615_5 gpc615_5_5402(
      {stage078[144], stage078[145], stage078[146], stage078[147], stage078[148]},
      {stage079[172]},
      {stage080[140], stage080[141], stage080[142], stage080[143], stage080[144], stage080[145]},
      {stage082[217], stage081[184], stage080[212], stage079[201], stage078[201]}
   );
   gpc615_5 gpc615_5_5403(
      {stage078[149], stage078[150], stage078[151], stage078[152], stage078[153]},
      {stage079[173]},
      {stage080[146], stage080[147], stage080[148], stage080[149], stage080[150], stage080[151]},
      {stage082[218], stage081[185], stage080[213], stage079[202], stage078[202]}
   );
   gpc615_5 gpc615_5_5404(
      {stage078[154], stage078[155], stage078[156], stage078[157], stage078[158]},
      {stage079[174]},
      {stage080[152], stage080[153], stage080[154], stage080[155], stage080[156], stage080[157]},
      {stage082[219], stage081[186], stage080[214], stage079[203], stage078[203]}
   );
   gpc615_5 gpc615_5_5405(
      {stage078[159], stage078[160], stage078[161], stage078[162], stage078[163]},
      {stage079[175]},
      {stage080[158], stage080[159], stage080[160], stage080[161], stage080[162], stage080[163]},
      {stage082[220], stage081[187], stage080[215], stage079[204], stage078[204]}
   );
   gpc615_5 gpc615_5_5406(
      {stage078[164], stage078[165], stage078[166], stage078[167], stage078[168]},
      {stage079[176]},
      {stage080[164], stage080[165], stage080[166], stage080[167], stage080[168], stage080[169]},
      {stage082[221], stage081[188], stage080[216], stage079[205], stage078[205]}
   );
   gpc615_5 gpc615_5_5407(
      {stage078[169], stage078[170], stage078[171], stage078[172], stage078[173]},
      {stage079[177]},
      {stage080[170], stage080[171], stage080[172], stage080[173], stage080[174], stage080[175]},
      {stage082[222], stage081[189], stage080[217], stage079[206], stage078[206]}
   );
   gpc1_1 gpc1_1_5408(
      {stage079[178]},
      {stage079[207]}
   );
   gpc1_1 gpc1_1_5409(
      {stage079[179]},
      {stage079[208]}
   );
   gpc1_1 gpc1_1_5410(
      {stage079[180]},
      {stage079[209]}
   );
   gpc1_1 gpc1_1_5411(
      {stage079[181]},
      {stage079[210]}
   );
   gpc1_1 gpc1_1_5412(
      {stage079[182]},
      {stage079[211]}
   );
   gpc1_1 gpc1_1_5413(
      {stage079[183]},
      {stage079[212]}
   );
   gpc1_1 gpc1_1_5414(
      {stage079[184]},
      {stage079[213]}
   );
   gpc1_1 gpc1_1_5415(
      {stage079[185]},
      {stage079[214]}
   );
   gpc1_1 gpc1_1_5416(
      {stage079[186]},
      {stage079[215]}
   );
   gpc1_1 gpc1_1_5417(
      {stage080[176]},
      {stage080[218]}
   );
   gpc1_1 gpc1_1_5418(
      {stage080[177]},
      {stage080[219]}
   );
   gpc1_1 gpc1_1_5419(
      {stage080[178]},
      {stage080[220]}
   );
   gpc1_1 gpc1_1_5420(
      {stage080[179]},
      {stage080[221]}
   );
   gpc1_1 gpc1_1_5421(
      {stage080[180]},
      {stage080[222]}
   );
   gpc1_1 gpc1_1_5422(
      {stage080[181]},
      {stage080[223]}
   );
   gpc1_1 gpc1_1_5423(
      {stage080[182]},
      {stage080[224]}
   );
   gpc1_1 gpc1_1_5424(
      {stage080[183]},
      {stage080[225]}
   );
   gpc1_1 gpc1_1_5425(
      {stage080[184]},
      {stage080[226]}
   );
   gpc1_1 gpc1_1_5426(
      {stage080[185]},
      {stage080[227]}
   );
   gpc1_1 gpc1_1_5427(
      {stage080[186]},
      {stage080[228]}
   );
   gpc606_5 gpc606_5_5428(
      {stage080[187], stage080[188], stage080[189], stage080[190], stage080[191], stage080[192]},
      {stage082[128], stage082[129], stage082[130], stage082[131], stage082[132], stage082[133]},
      {stage084[197], stage083[196], stage082[223], stage081[190], stage080[229]}
   );
   gpc615_5 gpc615_5_5429(
      {stage080[193], stage080[194], stage080[195], stage080[196], stage080[197]},
      {stage081[128]},
      {stage082[134], stage082[135], stage082[136], stage082[137], stage082[138], stage082[139]},
      {stage084[198], stage083[197], stage082[224], stage081[191], stage080[230]}
   );
   gpc615_5 gpc615_5_5430(
      {stage080[198], stage080[199], stage080[200], stage080[201], stage080[202]},
      {stage081[129]},
      {stage082[140], stage082[141], stage082[142], stage082[143], stage082[144], stage082[145]},
      {stage084[199], stage083[198], stage082[225], stage081[192], stage080[231]}
   );
   gpc1_1 gpc1_1_5431(
      {stage081[130]},
      {stage081[193]}
   );
   gpc1_1 gpc1_1_5432(
      {stage081[131]},
      {stage081[194]}
   );
   gpc1_1 gpc1_1_5433(
      {stage081[132]},
      {stage081[195]}
   );
   gpc1_1 gpc1_1_5434(
      {stage081[133]},
      {stage081[196]}
   );
   gpc1_1 gpc1_1_5435(
      {stage081[134]},
      {stage081[197]}
   );
   gpc1_1 gpc1_1_5436(
      {stage081[135]},
      {stage081[198]}
   );
   gpc1_1 gpc1_1_5437(
      {stage081[136]},
      {stage081[199]}
   );
   gpc1_1 gpc1_1_5438(
      {stage081[137]},
      {stage081[200]}
   );
   gpc1_1 gpc1_1_5439(
      {stage081[138]},
      {stage081[201]}
   );
   gpc1_1 gpc1_1_5440(
      {stage081[139]},
      {stage081[202]}
   );
   gpc1_1 gpc1_1_5441(
      {stage081[140]},
      {stage081[203]}
   );
   gpc1_1 gpc1_1_5442(
      {stage081[141]},
      {stage081[204]}
   );
   gpc1_1 gpc1_1_5443(
      {stage081[142]},
      {stage081[205]}
   );
   gpc1_1 gpc1_1_5444(
      {stage081[143]},
      {stage081[206]}
   );
   gpc1_1 gpc1_1_5445(
      {stage081[144]},
      {stage081[207]}
   );
   gpc1_1 gpc1_1_5446(
      {stage081[145]},
      {stage081[208]}
   );
   gpc1_1 gpc1_1_5447(
      {stage081[146]},
      {stage081[209]}
   );
   gpc1_1 gpc1_1_5448(
      {stage081[147]},
      {stage081[210]}
   );
   gpc1_1 gpc1_1_5449(
      {stage081[148]},
      {stage081[211]}
   );
   gpc1_1 gpc1_1_5450(
      {stage081[149]},
      {stage081[212]}
   );
   gpc1_1 gpc1_1_5451(
      {stage081[150]},
      {stage081[213]}
   );
   gpc1_1 gpc1_1_5452(
      {stage081[151]},
      {stage081[214]}
   );
   gpc1_1 gpc1_1_5453(
      {stage081[152]},
      {stage081[215]}
   );
   gpc1_1 gpc1_1_5454(
      {stage081[153]},
      {stage081[216]}
   );
   gpc1_1 gpc1_1_5455(
      {stage081[154]},
      {stage081[217]}
   );
   gpc1_1 gpc1_1_5456(
      {stage081[155]},
      {stage081[218]}
   );
   gpc1_1 gpc1_1_5457(
      {stage081[156]},
      {stage081[219]}
   );
   gpc1_1 gpc1_1_5458(
      {stage081[157]},
      {stage081[220]}
   );
   gpc1_1 gpc1_1_5459(
      {stage081[158]},
      {stage081[221]}
   );
   gpc1_1 gpc1_1_5460(
      {stage081[159]},
      {stage081[222]}
   );
   gpc1_1 gpc1_1_5461(
      {stage081[160]},
      {stage081[223]}
   );
   gpc1_1 gpc1_1_5462(
      {stage081[161]},
      {stage081[224]}
   );
   gpc1_1 gpc1_1_5463(
      {stage081[162]},
      {stage081[225]}
   );
   gpc1_1 gpc1_1_5464(
      {stage081[163]},
      {stage081[226]}
   );
   gpc1_1 gpc1_1_5465(
      {stage081[164]},
      {stage081[227]}
   );
   gpc1_1 gpc1_1_5466(
      {stage081[165]},
      {stage081[228]}
   );
   gpc1_1 gpc1_1_5467(
      {stage081[166]},
      {stage081[229]}
   );
   gpc1_1 gpc1_1_5468(
      {stage081[167]},
      {stage081[230]}
   );
   gpc1_1 gpc1_1_5469(
      {stage081[168]},
      {stage081[231]}
   );
   gpc1_1 gpc1_1_5470(
      {stage081[169]},
      {stage081[232]}
   );
   gpc1_1 gpc1_1_5471(
      {stage081[170]},
      {stage081[233]}
   );
   gpc1_1 gpc1_1_5472(
      {stage081[171]},
      {stage081[234]}
   );
   gpc1_1 gpc1_1_5473(
      {stage081[172]},
      {stage081[235]}
   );
   gpc1_1 gpc1_1_5474(
      {stage081[173]},
      {stage081[236]}
   );
   gpc1_1 gpc1_1_5475(
      {stage081[174]},
      {stage081[237]}
   );
   gpc1_1 gpc1_1_5476(
      {stage082[146]},
      {stage082[226]}
   );
   gpc1_1 gpc1_1_5477(
      {stage082[147]},
      {stage082[227]}
   );
   gpc1_1 gpc1_1_5478(
      {stage082[148]},
      {stage082[228]}
   );
   gpc606_5 gpc606_5_5479(
      {stage082[149], stage082[150], stage082[151], stage082[152], stage082[153], stage082[154]},
      {stage084[128], stage084[129], stage084[130], stage084[131], stage084[132], stage084[133]},
      {stage086[205], stage085[218], stage084[200], stage083[199], stage082[229]}
   );
   gpc606_5 gpc606_5_5480(
      {stage082[155], stage082[156], stage082[157], stage082[158], stage082[159], stage082[160]},
      {stage084[134], stage084[135], stage084[136], stage084[137], stage084[138], stage084[139]},
      {stage086[206], stage085[219], stage084[201], stage083[200], stage082[230]}
   );
   gpc606_5 gpc606_5_5481(
      {stage082[161], stage082[162], stage082[163], stage082[164], stage082[165], stage082[166]},
      {stage084[140], stage084[141], stage084[142], stage084[143], stage084[144], stage084[145]},
      {stage086[207], stage085[220], stage084[202], stage083[201], stage082[231]}
   );
   gpc606_5 gpc606_5_5482(
      {stage082[167], stage082[168], stage082[169], stage082[170], stage082[171], stage082[172]},
      {stage084[146], stage084[147], stage084[148], stage084[149], stage084[150], stage084[151]},
      {stage086[208], stage085[221], stage084[203], stage083[202], stage082[232]}
   );
   gpc606_5 gpc606_5_5483(
      {stage082[173], stage082[174], stage082[175], stage082[176], stage082[177], stage082[178]},
      {stage084[152], stage084[153], stage084[154], stage084[155], stage084[156], stage084[157]},
      {stage086[209], stage085[222], stage084[204], stage083[203], stage082[233]}
   );
   gpc606_5 gpc606_5_5484(
      {stage082[179], stage082[180], stage082[181], stage082[182], stage082[183], stage082[184]},
      {stage084[158], stage084[159], stage084[160], stage084[161], stage084[162], stage084[163]},
      {stage086[210], stage085[223], stage084[205], stage083[204], stage082[234]}
   );
   gpc606_5 gpc606_5_5485(
      {stage082[185], stage082[186], stage082[187], stage082[188], stage082[189], stage082[190]},
      {stage084[164], stage084[165], stage084[166], stage084[167], stage084[168], stage084[169]},
      {stage086[211], stage085[224], stage084[206], stage083[205], stage082[235]}
   );
   gpc606_5 gpc606_5_5486(
      {stage082[191], stage082[192], stage082[193], stage082[194], stage082[195], stage082[196]},
      {stage084[170], stage084[171], stage084[172], stage084[173], stage084[174], stage084[175]},
      {stage086[212], stage085[225], stage084[207], stage083[206], stage082[236]}
   );
   gpc606_5 gpc606_5_5487(
      {stage082[197], stage082[198], stage082[199], stage082[200], stage082[201], stage082[202]},
      {stage084[176], stage084[177], stage084[178], stage084[179], stage084[180], stage084[181]},
      {stage086[213], stage085[226], stage084[208], stage083[207], stage082[237]}
   );
   gpc606_5 gpc606_5_5488(
      {stage082[203], stage082[204], stage082[205], stage082[206], stage082[207], stage082[208]},
      {stage084[182], stage084[183], stage084[184], stage084[185], stage084[186], stage084[187]},
      {stage086[214], stage085[227], stage084[209], stage083[208], stage082[238]}
   );
   gpc606_5 gpc606_5_5489(
      {stage082[209], stage082[210], stage082[211], stage082[212], stage082[213], stage082[214]},
      {stage084[188], stage084[189], stage084[190], stage084[191], stage084[192], stage084[193]},
      {stage086[215], stage085[228], stage084[210], stage083[209], stage082[239]}
   );
   gpc1_1 gpc1_1_5490(
      {stage083[128]},
      {stage083[210]}
   );
   gpc1_1 gpc1_1_5491(
      {stage083[129]},
      {stage083[211]}
   );
   gpc1_1 gpc1_1_5492(
      {stage083[130]},
      {stage083[212]}
   );
   gpc1_1 gpc1_1_5493(
      {stage083[131]},
      {stage083[213]}
   );
   gpc1_1 gpc1_1_5494(
      {stage083[132]},
      {stage083[214]}
   );
   gpc1_1 gpc1_1_5495(
      {stage083[133]},
      {stage083[215]}
   );
   gpc1_1 gpc1_1_5496(
      {stage083[134]},
      {stage083[216]}
   );
   gpc1_1 gpc1_1_5497(
      {stage083[135]},
      {stage083[217]}
   );
   gpc1_1 gpc1_1_5498(
      {stage083[136]},
      {stage083[218]}
   );
   gpc1_1 gpc1_1_5499(
      {stage083[137]},
      {stage083[219]}
   );
   gpc1_1 gpc1_1_5500(
      {stage083[138]},
      {stage083[220]}
   );
   gpc1_1 gpc1_1_5501(
      {stage083[139]},
      {stage083[221]}
   );
   gpc1_1 gpc1_1_5502(
      {stage083[140]},
      {stage083[222]}
   );
   gpc1_1 gpc1_1_5503(
      {stage083[141]},
      {stage083[223]}
   );
   gpc1_1 gpc1_1_5504(
      {stage083[142]},
      {stage083[224]}
   );
   gpc1_1 gpc1_1_5505(
      {stage083[143]},
      {stage083[225]}
   );
   gpc1_1 gpc1_1_5506(
      {stage083[144]},
      {stage083[226]}
   );
   gpc1_1 gpc1_1_5507(
      {stage083[145]},
      {stage083[227]}
   );
   gpc1_1 gpc1_1_5508(
      {stage083[146]},
      {stage083[228]}
   );
   gpc1_1 gpc1_1_5509(
      {stage083[147]},
      {stage083[229]}
   );
   gpc1_1 gpc1_1_5510(
      {stage083[148]},
      {stage083[230]}
   );
   gpc1_1 gpc1_1_5511(
      {stage083[149]},
      {stage083[231]}
   );
   gpc1_1 gpc1_1_5512(
      {stage083[150]},
      {stage083[232]}
   );
   gpc1_1 gpc1_1_5513(
      {stage083[151]},
      {stage083[233]}
   );
   gpc1_1 gpc1_1_5514(
      {stage083[152]},
      {stage083[234]}
   );
   gpc1_1 gpc1_1_5515(
      {stage083[153]},
      {stage083[235]}
   );
   gpc1_1 gpc1_1_5516(
      {stage083[154]},
      {stage083[236]}
   );
   gpc1_1 gpc1_1_5517(
      {stage083[155]},
      {stage083[237]}
   );
   gpc1_1 gpc1_1_5518(
      {stage083[156]},
      {stage083[238]}
   );
   gpc606_5 gpc606_5_5519(
      {stage083[157], stage083[158], stage083[159], stage083[160], stage083[161], stage083[162]},
      {stage085[128], stage085[129], stage085[130], stage085[131], stage085[132], stage085[133]},
      {stage087[183], stage086[216], stage085[229], stage084[211], stage083[239]}
   );
   gpc606_5 gpc606_5_5520(
      {stage083[163], stage083[164], stage083[165], stage083[166], stage083[167], stage083[168]},
      {stage085[134], stage085[135], stage085[136], stage085[137], stage085[138], stage085[139]},
      {stage087[184], stage086[217], stage085[230], stage084[212], stage083[240]}
   );
   gpc606_5 gpc606_5_5521(
      {stage083[169], stage083[170], stage083[171], stage083[172], stage083[173], stage083[174]},
      {stage085[140], stage085[141], stage085[142], stage085[143], stage085[144], stage085[145]},
      {stage087[185], stage086[218], stage085[231], stage084[213], stage083[241]}
   );
   gpc606_5 gpc606_5_5522(
      {stage083[175], stage083[176], stage083[177], stage083[178], stage083[179], stage083[180]},
      {stage085[146], stage085[147], stage085[148], stage085[149], stage085[150], stage085[151]},
      {stage087[186], stage086[219], stage085[232], stage084[214], stage083[242]}
   );
   gpc615_5 gpc615_5_5523(
      {stage083[181], stage083[182], stage083[183], stage083[184], stage083[185]},
      {stage084[194]},
      {stage085[152], stage085[153], stage085[154], stage085[155], stage085[156], stage085[157]},
      {stage087[187], stage086[220], stage085[233], stage084[215], stage083[243]}
   );
   gpc615_5 gpc615_5_5524(
      {stage083[186], stage083[187], stage083[188], stage083[189], stage083[190]},
      {stage084[195]},
      {stage085[158], stage085[159], stage085[160], stage085[161], stage085[162], stage085[163]},
      {stage087[188], stage086[221], stage085[234], stage084[216], stage083[244]}
   );
   gpc615_5 gpc615_5_5525(
      {stage083[191], stage083[192], stage083[193], stage083[194], stage083[195]},
      {stage084[196]},
      {stage085[164], stage085[165], stage085[166], stage085[167], stage085[168], stage085[169]},
      {stage087[189], stage086[222], stage085[235], stage084[217], stage083[245]}
   );
   gpc1_1 gpc1_1_5526(
      {stage085[170]},
      {stage085[236]}
   );
   gpc1_1 gpc1_1_5527(
      {stage085[171]},
      {stage085[237]}
   );
   gpc1_1 gpc1_1_5528(
      {stage085[172]},
      {stage085[238]}
   );
   gpc1_1 gpc1_1_5529(
      {stage085[173]},
      {stage085[239]}
   );
   gpc1_1 gpc1_1_5530(
      {stage085[174]},
      {stage085[240]}
   );
   gpc1_1 gpc1_1_5531(
      {stage085[175]},
      {stage085[241]}
   );
   gpc606_5 gpc606_5_5532(
      {stage085[176], stage085[177], stage085[178], stage085[179], stage085[180], stage085[181]},
      {stage087[128], stage087[129], stage087[130], stage087[131], stage087[132], stage087[133]},
      {stage089[166], stage088[220], stage087[190], stage086[223], stage085[242]}
   );
   gpc606_5 gpc606_5_5533(
      {stage085[182], stage085[183], stage085[184], stage085[185], stage085[186], stage085[187]},
      {stage087[134], stage087[135], stage087[136], stage087[137], stage087[138], stage087[139]},
      {stage089[167], stage088[221], stage087[191], stage086[224], stage085[243]}
   );
   gpc606_5 gpc606_5_5534(
      {stage085[188], stage085[189], stage085[190], stage085[191], stage085[192], stage085[193]},
      {stage087[140], stage087[141], stage087[142], stage087[143], stage087[144], stage087[145]},
      {stage089[168], stage088[222], stage087[192], stage086[225], stage085[244]}
   );
   gpc606_5 gpc606_5_5535(
      {stage085[194], stage085[195], stage085[196], stage085[197], stage085[198], stage085[199]},
      {stage087[146], stage087[147], stage087[148], stage087[149], stage087[150], stage087[151]},
      {stage089[169], stage088[223], stage087[193], stage086[226], stage085[245]}
   );
   gpc606_5 gpc606_5_5536(
      {stage085[200], stage085[201], stage085[202], stage085[203], stage085[204], stage085[205]},
      {stage087[152], stage087[153], stage087[154], stage087[155], stage087[156], stage087[157]},
      {stage089[170], stage088[224], stage087[194], stage086[227], stage085[246]}
   );
   gpc606_5 gpc606_5_5537(
      {stage085[206], stage085[207], stage085[208], stage085[209], stage085[210], stage085[211]},
      {stage087[158], stage087[159], stage087[160], stage087[161], stage087[162], stage087[163]},
      {stage089[171], stage088[225], stage087[195], stage086[228], stage085[247]}
   );
   gpc606_5 gpc606_5_5538(
      {stage085[212], stage085[213], stage085[214], stage085[215], stage085[216], stage085[217]},
      {stage087[164], stage087[165], stage087[166], stage087[167], stage087[168], stage087[169]},
      {stage089[172], stage088[226], stage087[196], stage086[229], stage085[248]}
   );
   gpc606_5 gpc606_5_5539(
      {stage086[128], stage086[129], stage086[130], stage086[131], stage086[132], stage086[133]},
      {stage088[128], stage088[129], stage088[130], stage088[131], stage088[132], stage088[133]},
      {stage090[180], stage089[173], stage088[227], stage087[197], stage086[230]}
   );
   gpc606_5 gpc606_5_5540(
      {stage086[134], stage086[135], stage086[136], stage086[137], stage086[138], stage086[139]},
      {stage088[134], stage088[135], stage088[136], stage088[137], stage088[138], stage088[139]},
      {stage090[181], stage089[174], stage088[228], stage087[198], stage086[231]}
   );
   gpc606_5 gpc606_5_5541(
      {stage086[140], stage086[141], stage086[142], stage086[143], stage086[144], stage086[145]},
      {stage088[140], stage088[141], stage088[142], stage088[143], stage088[144], stage088[145]},
      {stage090[182], stage089[175], stage088[229], stage087[199], stage086[232]}
   );
   gpc606_5 gpc606_5_5542(
      {stage086[146], stage086[147], stage086[148], stage086[149], stage086[150], stage086[151]},
      {stage088[146], stage088[147], stage088[148], stage088[149], stage088[150], stage088[151]},
      {stage090[183], stage089[176], stage088[230], stage087[200], stage086[233]}
   );
   gpc606_5 gpc606_5_5543(
      {stage086[152], stage086[153], stage086[154], stage086[155], stage086[156], stage086[157]},
      {stage088[152], stage088[153], stage088[154], stage088[155], stage088[156], stage088[157]},
      {stage090[184], stage089[177], stage088[231], stage087[201], stage086[234]}
   );
   gpc606_5 gpc606_5_5544(
      {stage086[158], stage086[159], stage086[160], stage086[161], stage086[162], stage086[163]},
      {stage088[158], stage088[159], stage088[160], stage088[161], stage088[162], stage088[163]},
      {stage090[185], stage089[178], stage088[232], stage087[202], stage086[235]}
   );
   gpc606_5 gpc606_5_5545(
      {stage086[164], stage086[165], stage086[166], stage086[167], stage086[168], stage086[169]},
      {stage088[164], stage088[165], stage088[166], stage088[167], stage088[168], stage088[169]},
      {stage090[186], stage089[179], stage088[233], stage087[203], stage086[236]}
   );
   gpc606_5 gpc606_5_5546(
      {stage086[170], stage086[171], stage086[172], stage086[173], stage086[174], stage086[175]},
      {stage088[170], stage088[171], stage088[172], stage088[173], stage088[174], stage088[175]},
      {stage090[187], stage089[180], stage088[234], stage087[204], stage086[237]}
   );
   gpc606_5 gpc606_5_5547(
      {stage086[176], stage086[177], stage086[178], stage086[179], stage086[180], stage086[181]},
      {stage088[176], stage088[177], stage088[178], stage088[179], stage088[180], stage088[181]},
      {stage090[188], stage089[181], stage088[235], stage087[205], stage086[238]}
   );
   gpc606_5 gpc606_5_5548(
      {stage086[182], stage086[183], stage086[184], stage086[185], stage086[186], stage086[187]},
      {stage088[182], stage088[183], stage088[184], stage088[185], stage088[186], stage088[187]},
      {stage090[189], stage089[182], stage088[236], stage087[206], stage086[239]}
   );
   gpc606_5 gpc606_5_5549(
      {stage086[188], stage086[189], stage086[190], stage086[191], stage086[192], stage086[193]},
      {stage088[188], stage088[189], stage088[190], stage088[191], stage088[192], stage088[193]},
      {stage090[190], stage089[183], stage088[237], stage087[207], stage086[240]}
   );
   gpc606_5 gpc606_5_5550(
      {stage086[194], stage086[195], stage086[196], stage086[197], stage086[198], stage086[199]},
      {stage088[194], stage088[195], stage088[196], stage088[197], stage088[198], stage088[199]},
      {stage090[191], stage089[184], stage088[238], stage087[208], stage086[241]}
   );
   gpc606_5 gpc606_5_5551(
      {stage086[200], stage086[201], stage086[202], stage086[203], stage086[204], 1'h0},
      {stage088[200], stage088[201], stage088[202], stage088[203], stage088[204], stage088[205]},
      {stage090[192], stage089[185], stage088[239], stage087[209], stage086[242]}
   );
   gpc1_1 gpc1_1_5552(
      {stage087[170]},
      {stage087[210]}
   );
   gpc606_5 gpc606_5_5553(
      {stage087[171], stage087[172], stage087[173], stage087[174], stage087[175], stage087[176]},
      {stage089[128], stage089[129], stage089[130], stage089[131], stage089[132], stage089[133]},
      {stage091[200], stage090[193], stage089[186], stage088[240], stage087[211]}
   );
   gpc606_5 gpc606_5_5554(
      {stage087[177], stage087[178], stage087[179], stage087[180], stage087[181], stage087[182]},
      {stage089[134], stage089[135], stage089[136], stage089[137], stage089[138], stage089[139]},
      {stage091[201], stage090[194], stage089[187], stage088[241], stage087[212]}
   );
   gpc1_1 gpc1_1_5555(
      {stage088[206]},
      {stage088[242]}
   );
   gpc1_1 gpc1_1_5556(
      {stage088[207]},
      {stage088[243]}
   );
   gpc606_5 gpc606_5_5557(
      {stage088[208], stage088[209], stage088[210], stage088[211], stage088[212], stage088[213]},
      {stage090[128], stage090[129], stage090[130], stage090[131], stage090[132], stage090[133]},
      {stage092[198], stage091[202], stage090[195], stage089[188], stage088[244]}
   );
   gpc606_5 gpc606_5_5558(
      {stage088[214], stage088[215], stage088[216], stage088[217], stage088[218], stage088[219]},
      {stage090[134], stage090[135], stage090[136], stage090[137], stage090[138], stage090[139]},
      {stage092[199], stage091[203], stage090[196], stage089[189], stage088[245]}
   );
   gpc1_1 gpc1_1_5559(
      {stage089[140]},
      {stage089[190]}
   );
   gpc1_1 gpc1_1_5560(
      {stage089[141]},
      {stage089[191]}
   );
   gpc1_1 gpc1_1_5561(
      {stage089[142]},
      {stage089[192]}
   );
   gpc1_1 gpc1_1_5562(
      {stage089[143]},
      {stage089[193]}
   );
   gpc1_1 gpc1_1_5563(
      {stage089[144]},
      {stage089[194]}
   );
   gpc1_1 gpc1_1_5564(
      {stage089[145]},
      {stage089[195]}
   );
   gpc1_1 gpc1_1_5565(
      {stage089[146]},
      {stage089[196]}
   );
   gpc1_1 gpc1_1_5566(
      {stage089[147]},
      {stage089[197]}
   );
   gpc1_1 gpc1_1_5567(
      {stage089[148]},
      {stage089[198]}
   );
   gpc1_1 gpc1_1_5568(
      {stage089[149]},
      {stage089[199]}
   );
   gpc1_1 gpc1_1_5569(
      {stage089[150]},
      {stage089[200]}
   );
   gpc1_1 gpc1_1_5570(
      {stage089[151]},
      {stage089[201]}
   );
   gpc1_1 gpc1_1_5571(
      {stage089[152]},
      {stage089[202]}
   );
   gpc1_1 gpc1_1_5572(
      {stage089[153]},
      {stage089[203]}
   );
   gpc1_1 gpc1_1_5573(
      {stage089[154]},
      {stage089[204]}
   );
   gpc1_1 gpc1_1_5574(
      {stage089[155]},
      {stage089[205]}
   );
   gpc1_1 gpc1_1_5575(
      {stage089[156]},
      {stage089[206]}
   );
   gpc1_1 gpc1_1_5576(
      {stage089[157]},
      {stage089[207]}
   );
   gpc1_1 gpc1_1_5577(
      {stage089[158]},
      {stage089[208]}
   );
   gpc1_1 gpc1_1_5578(
      {stage089[159]},
      {stage089[209]}
   );
   gpc1_1 gpc1_1_5579(
      {stage089[160]},
      {stage089[210]}
   );
   gpc1_1 gpc1_1_5580(
      {stage089[161]},
      {stage089[211]}
   );
   gpc1_1 gpc1_1_5581(
      {stage089[162]},
      {stage089[212]}
   );
   gpc1_1 gpc1_1_5582(
      {stage089[163]},
      {stage089[213]}
   );
   gpc1_1 gpc1_1_5583(
      {stage089[164]},
      {stage089[214]}
   );
   gpc1_1 gpc1_1_5584(
      {stage089[165]},
      {stage089[215]}
   );
   gpc1_1 gpc1_1_5585(
      {stage090[140]},
      {stage090[197]}
   );
   gpc1_1 gpc1_1_5586(
      {stage090[141]},
      {stage090[198]}
   );
   gpc1_1 gpc1_1_5587(
      {stage090[142]},
      {stage090[199]}
   );
   gpc1_1 gpc1_1_5588(
      {stage090[143]},
      {stage090[200]}
   );
   gpc1_1 gpc1_1_5589(
      {stage090[144]},
      {stage090[201]}
   );
   gpc1_1 gpc1_1_5590(
      {stage090[145]},
      {stage090[202]}
   );
   gpc1_1 gpc1_1_5591(
      {stage090[146]},
      {stage090[203]}
   );
   gpc1_1 gpc1_1_5592(
      {stage090[147]},
      {stage090[204]}
   );
   gpc1_1 gpc1_1_5593(
      {stage090[148]},
      {stage090[205]}
   );
   gpc1_1 gpc1_1_5594(
      {stage090[149]},
      {stage090[206]}
   );
   gpc1_1 gpc1_1_5595(
      {stage090[150]},
      {stage090[207]}
   );
   gpc1_1 gpc1_1_5596(
      {stage090[151]},
      {stage090[208]}
   );
   gpc1_1 gpc1_1_5597(
      {stage090[152]},
      {stage090[209]}
   );
   gpc1_1 gpc1_1_5598(
      {stage090[153]},
      {stage090[210]}
   );
   gpc1_1 gpc1_1_5599(
      {stage090[154]},
      {stage090[211]}
   );
   gpc1_1 gpc1_1_5600(
      {stage090[155]},
      {stage090[212]}
   );
   gpc606_5 gpc606_5_5601(
      {stage090[156], stage090[157], stage090[158], stage090[159], stage090[160], stage090[161]},
      {stage092[128], stage092[129], stage092[130], stage092[131], stage092[132], stage092[133]},
      {stage094[195], stage093[189], stage092[200], stage091[204], stage090[213]}
   );
   gpc606_5 gpc606_5_5602(
      {stage090[162], stage090[163], stage090[164], stage090[165], stage090[166], stage090[167]},
      {stage092[134], stage092[135], stage092[136], stage092[137], stage092[138], stage092[139]},
      {stage094[196], stage093[190], stage092[201], stage091[205], stage090[214]}
   );
   gpc606_5 gpc606_5_5603(
      {stage090[168], stage090[169], stage090[170], stage090[171], stage090[172], stage090[173]},
      {stage092[140], stage092[141], stage092[142], stage092[143], stage092[144], stage092[145]},
      {stage094[197], stage093[191], stage092[202], stage091[206], stage090[215]}
   );
   gpc606_5 gpc606_5_5604(
      {stage090[174], stage090[175], stage090[176], stage090[177], stage090[178], stage090[179]},
      {stage092[146], stage092[147], stage092[148], stage092[149], stage092[150], stage092[151]},
      {stage094[198], stage093[192], stage092[203], stage091[207], stage090[216]}
   );
   gpc1_1 gpc1_1_5605(
      {stage091[128]},
      {stage091[208]}
   );
   gpc1_1 gpc1_1_5606(
      {stage091[129]},
      {stage091[209]}
   );
   gpc1_1 gpc1_1_5607(
      {stage091[130]},
      {stage091[210]}
   );
   gpc1_1 gpc1_1_5608(
      {stage091[131]},
      {stage091[211]}
   );
   gpc1_1 gpc1_1_5609(
      {stage091[132]},
      {stage091[212]}
   );
   gpc1_1 gpc1_1_5610(
      {stage091[133]},
      {stage091[213]}
   );
   gpc1_1 gpc1_1_5611(
      {stage091[134]},
      {stage091[214]}
   );
   gpc1_1 gpc1_1_5612(
      {stage091[135]},
      {stage091[215]}
   );
   gpc1_1 gpc1_1_5613(
      {stage091[136]},
      {stage091[216]}
   );
   gpc1_1 gpc1_1_5614(
      {stage091[137]},
      {stage091[217]}
   );
   gpc1_1 gpc1_1_5615(
      {stage091[138]},
      {stage091[218]}
   );
   gpc1_1 gpc1_1_5616(
      {stage091[139]},
      {stage091[219]}
   );
   gpc1_1 gpc1_1_5617(
      {stage091[140]},
      {stage091[220]}
   );
   gpc1_1 gpc1_1_5618(
      {stage091[141]},
      {stage091[221]}
   );
   gpc1_1 gpc1_1_5619(
      {stage091[142]},
      {stage091[222]}
   );
   gpc1_1 gpc1_1_5620(
      {stage091[143]},
      {stage091[223]}
   );
   gpc1_1 gpc1_1_5621(
      {stage091[144]},
      {stage091[224]}
   );
   gpc1_1 gpc1_1_5622(
      {stage091[145]},
      {stage091[225]}
   );
   gpc1_1 gpc1_1_5623(
      {stage091[146]},
      {stage091[226]}
   );
   gpc1_1 gpc1_1_5624(
      {stage091[147]},
      {stage091[227]}
   );
   gpc1_1 gpc1_1_5625(
      {stage091[148]},
      {stage091[228]}
   );
   gpc1_1 gpc1_1_5626(
      {stage091[149]},
      {stage091[229]}
   );
   gpc1_1 gpc1_1_5627(
      {stage091[150]},
      {stage091[230]}
   );
   gpc1_1 gpc1_1_5628(
      {stage091[151]},
      {stage091[231]}
   );
   gpc1_1 gpc1_1_5629(
      {stage091[152]},
      {stage091[232]}
   );
   gpc1_1 gpc1_1_5630(
      {stage091[153]},
      {stage091[233]}
   );
   gpc1_1 gpc1_1_5631(
      {stage091[154]},
      {stage091[234]}
   );
   gpc1_1 gpc1_1_5632(
      {stage091[155]},
      {stage091[235]}
   );
   gpc1_1 gpc1_1_5633(
      {stage091[156]},
      {stage091[236]}
   );
   gpc1_1 gpc1_1_5634(
      {stage091[157]},
      {stage091[237]}
   );
   gpc1_1 gpc1_1_5635(
      {stage091[158]},
      {stage091[238]}
   );
   gpc1_1 gpc1_1_5636(
      {stage091[159]},
      {stage091[239]}
   );
   gpc1_1 gpc1_1_5637(
      {stage091[160]},
      {stage091[240]}
   );
   gpc1_1 gpc1_1_5638(
      {stage091[161]},
      {stage091[241]}
   );
   gpc1_1 gpc1_1_5639(
      {stage091[162]},
      {stage091[242]}
   );
   gpc1_1 gpc1_1_5640(
      {stage091[163]},
      {stage091[243]}
   );
   gpc1_1 gpc1_1_5641(
      {stage091[164]},
      {stage091[244]}
   );
   gpc1_1 gpc1_1_5642(
      {stage091[165]},
      {stage091[245]}
   );
   gpc1_1 gpc1_1_5643(
      {stage091[166]},
      {stage091[246]}
   );
   gpc1_1 gpc1_1_5644(
      {stage091[167]},
      {stage091[247]}
   );
   gpc1_1 gpc1_1_5645(
      {stage091[168]},
      {stage091[248]}
   );
   gpc1_1 gpc1_1_5646(
      {stage091[169]},
      {stage091[249]}
   );
   gpc606_5 gpc606_5_5647(
      {stage091[170], stage091[171], stage091[172], stage091[173], stage091[174], stage091[175]},
      {stage093[128], stage093[129], stage093[130], stage093[131], stage093[132], stage093[133]},
      {stage095[181], stage094[199], stage093[193], stage092[204], stage091[250]}
   );
   gpc606_5 gpc606_5_5648(
      {stage091[176], stage091[177], stage091[178], stage091[179], stage091[180], stage091[181]},
      {stage093[134], stage093[135], stage093[136], stage093[137], stage093[138], stage093[139]},
      {stage095[182], stage094[200], stage093[194], stage092[205], stage091[251]}
   );
   gpc606_5 gpc606_5_5649(
      {stage091[182], stage091[183], stage091[184], stage091[185], stage091[186], stage091[187]},
      {stage093[140], stage093[141], stage093[142], stage093[143], stage093[144], stage093[145]},
      {stage095[183], stage094[201], stage093[195], stage092[206], stage091[252]}
   );
   gpc606_5 gpc606_5_5650(
      {stage091[188], stage091[189], stage091[190], stage091[191], stage091[192], stage091[193]},
      {stage093[146], stage093[147], stage093[148], stage093[149], stage093[150], stage093[151]},
      {stage095[184], stage094[202], stage093[196], stage092[207], stage091[253]}
   );
   gpc606_5 gpc606_5_5651(
      {stage091[194], stage091[195], stage091[196], stage091[197], stage091[198], stage091[199]},
      {stage093[152], stage093[153], stage093[154], stage093[155], stage093[156], stage093[157]},
      {stage095[185], stage094[203], stage093[197], stage092[208], stage091[254]}
   );
   gpc1_1 gpc1_1_5652(
      {stage092[152]},
      {stage092[209]}
   );
   gpc1_1 gpc1_1_5653(
      {stage092[153]},
      {stage092[210]}
   );
   gpc1_1 gpc1_1_5654(
      {stage092[154]},
      {stage092[211]}
   );
   gpc1_1 gpc1_1_5655(
      {stage092[155]},
      {stage092[212]}
   );
   gpc1_1 gpc1_1_5656(
      {stage092[156]},
      {stage092[213]}
   );
   gpc1_1 gpc1_1_5657(
      {stage092[157]},
      {stage092[214]}
   );
   gpc1_1 gpc1_1_5658(
      {stage092[158]},
      {stage092[215]}
   );
   gpc1_1 gpc1_1_5659(
      {stage092[159]},
      {stage092[216]}
   );
   gpc1_1 gpc1_1_5660(
      {stage092[160]},
      {stage092[217]}
   );
   gpc1_1 gpc1_1_5661(
      {stage092[161]},
      {stage092[218]}
   );
   gpc1_1 gpc1_1_5662(
      {stage092[162]},
      {stage092[219]}
   );
   gpc615_5 gpc615_5_5663(
      {stage092[163], stage092[164], stage092[165], stage092[166], stage092[167]},
      {stage093[158]},
      {stage094[128], stage094[129], stage094[130], stage094[131], stage094[132], stage094[133]},
      {stage096[184], stage095[186], stage094[204], stage093[198], stage092[220]}
   );
   gpc615_5 gpc615_5_5664(
      {stage092[168], stage092[169], stage092[170], stage092[171], stage092[172]},
      {stage093[159]},
      {stage094[134], stage094[135], stage094[136], stage094[137], stage094[138], stage094[139]},
      {stage096[185], stage095[187], stage094[205], stage093[199], stage092[221]}
   );
   gpc615_5 gpc615_5_5665(
      {stage092[173], stage092[174], stage092[175], stage092[176], stage092[177]},
      {stage093[160]},
      {stage094[140], stage094[141], stage094[142], stage094[143], stage094[144], stage094[145]},
      {stage096[186], stage095[188], stage094[206], stage093[200], stage092[222]}
   );
   gpc615_5 gpc615_5_5666(
      {stage092[178], stage092[179], stage092[180], stage092[181], stage092[182]},
      {stage093[161]},
      {stage094[146], stage094[147], stage094[148], stage094[149], stage094[150], stage094[151]},
      {stage096[187], stage095[189], stage094[207], stage093[201], stage092[223]}
   );
   gpc615_5 gpc615_5_5667(
      {stage092[183], stage092[184], stage092[185], stage092[186], stage092[187]},
      {stage093[162]},
      {stage094[152], stage094[153], stage094[154], stage094[155], stage094[156], stage094[157]},
      {stage096[188], stage095[190], stage094[208], stage093[202], stage092[224]}
   );
   gpc615_5 gpc615_5_5668(
      {stage092[188], stage092[189], stage092[190], stage092[191], stage092[192]},
      {stage093[163]},
      {stage094[158], stage094[159], stage094[160], stage094[161], stage094[162], stage094[163]},
      {stage096[189], stage095[191], stage094[209], stage093[203], stage092[225]}
   );
   gpc615_5 gpc615_5_5669(
      {stage092[193], stage092[194], stage092[195], stage092[196], stage092[197]},
      {stage093[164]},
      {stage094[164], stage094[165], stage094[166], stage094[167], stage094[168], stage094[169]},
      {stage096[190], stage095[192], stage094[210], stage093[204], stage092[226]}
   );
   gpc606_5 gpc606_5_5670(
      {stage093[165], stage093[166], stage093[167], stage093[168], stage093[169], stage093[170]},
      {stage095[128], stage095[129], stage095[130], stage095[131], stage095[132], stage095[133]},
      {stage097[175], stage096[191], stage095[193], stage094[211], stage093[205]}
   );
   gpc606_5 gpc606_5_5671(
      {stage093[171], stage093[172], stage093[173], stage093[174], stage093[175], stage093[176]},
      {stage095[134], stage095[135], stage095[136], stage095[137], stage095[138], stage095[139]},
      {stage097[176], stage096[192], stage095[194], stage094[212], stage093[206]}
   );
   gpc606_5 gpc606_5_5672(
      {stage093[177], stage093[178], stage093[179], stage093[180], stage093[181], stage093[182]},
      {stage095[140], stage095[141], stage095[142], stage095[143], stage095[144], stage095[145]},
      {stage097[177], stage096[193], stage095[195], stage094[213], stage093[207]}
   );
   gpc606_5 gpc606_5_5673(
      {stage093[183], stage093[184], stage093[185], stage093[186], stage093[187], stage093[188]},
      {stage095[146], stage095[147], stage095[148], stage095[149], stage095[150], stage095[151]},
      {stage097[178], stage096[194], stage095[196], stage094[214], stage093[208]}
   );
   gpc1_1 gpc1_1_5674(
      {stage094[170]},
      {stage094[215]}
   );
   gpc1_1 gpc1_1_5675(
      {stage094[171]},
      {stage094[216]}
   );
   gpc1_1 gpc1_1_5676(
      {stage094[172]},
      {stage094[217]}
   );
   gpc1_1 gpc1_1_5677(
      {stage094[173]},
      {stage094[218]}
   );
   gpc1_1 gpc1_1_5678(
      {stage094[174]},
      {stage094[219]}
   );
   gpc1_1 gpc1_1_5679(
      {stage094[175]},
      {stage094[220]}
   );
   gpc7_3 gpc7_3_5680(
      {stage094[176], stage094[177], stage094[178], stage094[179], stage094[180], stage094[181], stage094[182]},
      {stage096[195], stage095[197], stage094[221]}
   );
   gpc606_5 gpc606_5_5681(
      {stage094[183], stage094[184], stage094[185], stage094[186], stage094[187], stage094[188]},
      {stage096[128], stage096[129], stage096[130], stage096[131], stage096[132], stage096[133]},
      {stage098[184], stage097[179], stage096[196], stage095[198], stage094[222]}
   );
   gpc606_5 gpc606_5_5682(
      {stage094[189], stage094[190], stage094[191], stage094[192], stage094[193], stage094[194]},
      {stage096[134], stage096[135], stage096[136], stage096[137], stage096[138], stage096[139]},
      {stage098[185], stage097[180], stage096[197], stage095[199], stage094[223]}
   );
   gpc606_5 gpc606_5_5683(
      {stage095[152], stage095[153], stage095[154], stage095[155], stage095[156], stage095[157]},
      {stage097[128], stage097[129], stage097[130], stage097[131], stage097[132], stage097[133]},
      {stage099[204], stage098[186], stage097[181], stage096[198], stage095[200]}
   );
   gpc606_5 gpc606_5_5684(
      {stage095[158], stage095[159], stage095[160], stage095[161], stage095[162], stage095[163]},
      {stage097[134], stage097[135], stage097[136], stage097[137], stage097[138], stage097[139]},
      {stage099[205], stage098[187], stage097[182], stage096[199], stage095[201]}
   );
   gpc606_5 gpc606_5_5685(
      {stage095[164], stage095[165], stage095[166], stage095[167], stage095[168], stage095[169]},
      {stage097[140], stage097[141], stage097[142], stage097[143], stage097[144], stage097[145]},
      {stage099[206], stage098[188], stage097[183], stage096[200], stage095[202]}
   );
   gpc606_5 gpc606_5_5686(
      {stage095[170], stage095[171], stage095[172], stage095[173], stage095[174], stage095[175]},
      {stage097[146], stage097[147], stage097[148], stage097[149], stage097[150], stage097[151]},
      {stage099[207], stage098[189], stage097[184], stage096[201], stage095[203]}
   );
   gpc1415_5 gpc1415_5_5687(
      {stage095[176], stage095[177], stage095[178], stage095[179], stage095[180]},
      {stage096[140]},
      {stage097[152], stage097[153], stage097[154], stage097[155]},
      {stage098[128]},
      {stage099[208], stage098[190], stage097[185], stage096[202], stage095[204]}
   );
   gpc1_1 gpc1_1_5688(
      {stage096[141]},
      {stage096[203]}
   );
   gpc1_1 gpc1_1_5689(
      {stage096[142]},
      {stage096[204]}
   );
   gpc1_1 gpc1_1_5690(
      {stage096[143]},
      {stage096[205]}
   );
   gpc1_1 gpc1_1_5691(
      {stage096[144]},
      {stage096[206]}
   );
   gpc1_1 gpc1_1_5692(
      {stage096[145]},
      {stage096[207]}
   );
   gpc1_1 gpc1_1_5693(
      {stage096[146]},
      {stage096[208]}
   );
   gpc1_1 gpc1_1_5694(
      {stage096[147]},
      {stage096[209]}
   );
   gpc1_1 gpc1_1_5695(
      {stage096[148]},
      {stage096[210]}
   );
   gpc615_5 gpc615_5_5696(
      {stage096[149], stage096[150], stage096[151], stage096[152], stage096[153]},
      {stage097[156]},
      {stage098[129], stage098[130], stage098[131], stage098[132], stage098[133], stage098[134]},
      {stage100[178], stage099[209], stage098[191], stage097[186], stage096[211]}
   );
   gpc615_5 gpc615_5_5697(
      {stage096[154], stage096[155], stage096[156], stage096[157], stage096[158]},
      {stage097[157]},
      {stage098[135], stage098[136], stage098[137], stage098[138], stage098[139], stage098[140]},
      {stage100[179], stage099[210], stage098[192], stage097[187], stage096[212]}
   );
   gpc615_5 gpc615_5_5698(
      {stage096[159], stage096[160], stage096[161], stage096[162], stage096[163]},
      {stage097[158]},
      {stage098[141], stage098[142], stage098[143], stage098[144], stage098[145], stage098[146]},
      {stage100[180], stage099[211], stage098[193], stage097[188], stage096[213]}
   );
   gpc615_5 gpc615_5_5699(
      {stage096[164], stage096[165], stage096[166], stage096[167], stage096[168]},
      {stage097[159]},
      {stage098[147], stage098[148], stage098[149], stage098[150], stage098[151], stage098[152]},
      {stage100[181], stage099[212], stage098[194], stage097[189], stage096[214]}
   );
   gpc615_5 gpc615_5_5700(
      {stage096[169], stage096[170], stage096[171], stage096[172], stage096[173]},
      {stage097[160]},
      {stage098[153], stage098[154], stage098[155], stage098[156], stage098[157], stage098[158]},
      {stage100[182], stage099[213], stage098[195], stage097[190], stage096[215]}
   );
   gpc615_5 gpc615_5_5701(
      {stage096[174], stage096[175], stage096[176], stage096[177], stage096[178]},
      {stage097[161]},
      {stage098[159], stage098[160], stage098[161], stage098[162], stage098[163], stage098[164]},
      {stage100[183], stage099[214], stage098[196], stage097[191], stage096[216]}
   );
   gpc615_5 gpc615_5_5702(
      {stage096[179], stage096[180], stage096[181], stage096[182], stage096[183]},
      {stage097[162]},
      {stage098[165], stage098[166], stage098[167], stage098[168], stage098[169], stage098[170]},
      {stage100[184], stage099[215], stage098[197], stage097[192], stage096[217]}
   );
   gpc1_1 gpc1_1_5703(
      {stage097[163]},
      {stage097[193]}
   );
   gpc1_1 gpc1_1_5704(
      {stage097[164]},
      {stage097[194]}
   );
   gpc1_1 gpc1_1_5705(
      {stage097[165]},
      {stage097[195]}
   );
   gpc1_1 gpc1_1_5706(
      {stage097[166]},
      {stage097[196]}
   );
   gpc1_1 gpc1_1_5707(
      {stage097[167]},
      {stage097[197]}
   );
   gpc1_1 gpc1_1_5708(
      {stage097[168]},
      {stage097[198]}
   );
   gpc1_1 gpc1_1_5709(
      {stage097[169]},
      {stage097[199]}
   );
   gpc1_1 gpc1_1_5710(
      {stage097[170]},
      {stage097[200]}
   );
   gpc1_1 gpc1_1_5711(
      {stage097[171]},
      {stage097[201]}
   );
   gpc1_1 gpc1_1_5712(
      {stage097[172]},
      {stage097[202]}
   );
   gpc1_1 gpc1_1_5713(
      {stage097[173]},
      {stage097[203]}
   );
   gpc1_1 gpc1_1_5714(
      {stage097[174]},
      {stage097[204]}
   );
   gpc1_1 gpc1_1_5715(
      {stage098[171]},
      {stage098[198]}
   );
   gpc1_1 gpc1_1_5716(
      {stage098[172]},
      {stage098[199]}
   );
   gpc1_1 gpc1_1_5717(
      {stage098[173]},
      {stage098[200]}
   );
   gpc1_1 gpc1_1_5718(
      {stage098[174]},
      {stage098[201]}
   );
   gpc1_1 gpc1_1_5719(
      {stage098[175]},
      {stage098[202]}
   );
   gpc1_1 gpc1_1_5720(
      {stage098[176]},
      {stage098[203]}
   );
   gpc1_1 gpc1_1_5721(
      {stage098[177]},
      {stage098[204]}
   );
   gpc606_5 gpc606_5_5722(
      {stage098[178], stage098[179], stage098[180], stage098[181], stage098[182], stage098[183]},
      {stage100[128], stage100[129], stage100[130], stage100[131], stage100[132], stage100[133]},
      {stage102[200], stage101[192], stage100[185], stage099[216], stage098[205]}
   );
   gpc1_1 gpc1_1_5723(
      {stage099[128]},
      {stage099[217]}
   );
   gpc1_1 gpc1_1_5724(
      {stage099[129]},
      {stage099[218]}
   );
   gpc1_1 gpc1_1_5725(
      {stage099[130]},
      {stage099[219]}
   );
   gpc1_1 gpc1_1_5726(
      {stage099[131]},
      {stage099[220]}
   );
   gpc1_1 gpc1_1_5727(
      {stage099[132]},
      {stage099[221]}
   );
   gpc1_1 gpc1_1_5728(
      {stage099[133]},
      {stage099[222]}
   );
   gpc1_1 gpc1_1_5729(
      {stage099[134]},
      {stage099[223]}
   );
   gpc1_1 gpc1_1_5730(
      {stage099[135]},
      {stage099[224]}
   );
   gpc1_1 gpc1_1_5731(
      {stage099[136]},
      {stage099[225]}
   );
   gpc1_1 gpc1_1_5732(
      {stage099[137]},
      {stage099[226]}
   );
   gpc1_1 gpc1_1_5733(
      {stage099[138]},
      {stage099[227]}
   );
   gpc1_1 gpc1_1_5734(
      {stage099[139]},
      {stage099[228]}
   );
   gpc1_1 gpc1_1_5735(
      {stage099[140]},
      {stage099[229]}
   );
   gpc1_1 gpc1_1_5736(
      {stage099[141]},
      {stage099[230]}
   );
   gpc1_1 gpc1_1_5737(
      {stage099[142]},
      {stage099[231]}
   );
   gpc1_1 gpc1_1_5738(
      {stage099[143]},
      {stage099[232]}
   );
   gpc1_1 gpc1_1_5739(
      {stage099[144]},
      {stage099[233]}
   );
   gpc1_1 gpc1_1_5740(
      {stage099[145]},
      {stage099[234]}
   );
   gpc1_1 gpc1_1_5741(
      {stage099[146]},
      {stage099[235]}
   );
   gpc1_1 gpc1_1_5742(
      {stage099[147]},
      {stage099[236]}
   );
   gpc1_1 gpc1_1_5743(
      {stage099[148]},
      {stage099[237]}
   );
   gpc1_1 gpc1_1_5744(
      {stage099[149]},
      {stage099[238]}
   );
   gpc1_1 gpc1_1_5745(
      {stage099[150]},
      {stage099[239]}
   );
   gpc1_1 gpc1_1_5746(
      {stage099[151]},
      {stage099[240]}
   );
   gpc1_1 gpc1_1_5747(
      {stage099[152]},
      {stage099[241]}
   );
   gpc1_1 gpc1_1_5748(
      {stage099[153]},
      {stage099[242]}
   );
   gpc1_1 gpc1_1_5749(
      {stage099[154]},
      {stage099[243]}
   );
   gpc1_1 gpc1_1_5750(
      {stage099[155]},
      {stage099[244]}
   );
   gpc1_1 gpc1_1_5751(
      {stage099[156]},
      {stage099[245]}
   );
   gpc1_1 gpc1_1_5752(
      {stage099[157]},
      {stage099[246]}
   );
   gpc1_1 gpc1_1_5753(
      {stage099[158]},
      {stage099[247]}
   );
   gpc1_1 gpc1_1_5754(
      {stage099[159]},
      {stage099[248]}
   );
   gpc1_1 gpc1_1_5755(
      {stage099[160]},
      {stage099[249]}
   );
   gpc1_1 gpc1_1_5756(
      {stage099[161]},
      {stage099[250]}
   );
   gpc606_5 gpc606_5_5757(
      {stage099[162], stage099[163], stage099[164], stage099[165], stage099[166], stage099[167]},
      {stage101[128], stage101[129], stage101[130], stage101[131], stage101[132], stage101[133]},
      {stage103[192], stage102[201], stage101[193], stage100[186], stage099[251]}
   );
   gpc606_5 gpc606_5_5758(
      {stage099[168], stage099[169], stage099[170], stage099[171], stage099[172], stage099[173]},
      {stage101[134], stage101[135], stage101[136], stage101[137], stage101[138], stage101[139]},
      {stage103[193], stage102[202], stage101[194], stage100[187], stage099[252]}
   );
   gpc606_5 gpc606_5_5759(
      {stage099[174], stage099[175], stage099[176], stage099[177], stage099[178], stage099[179]},
      {stage101[140], stage101[141], stage101[142], stage101[143], stage101[144], stage101[145]},
      {stage103[194], stage102[203], stage101[195], stage100[188], stage099[253]}
   );
   gpc606_5 gpc606_5_5760(
      {stage099[180], stage099[181], stage099[182], stage099[183], stage099[184], stage099[185]},
      {stage101[146], stage101[147], stage101[148], stage101[149], stage101[150], stage101[151]},
      {stage103[195], stage102[204], stage101[196], stage100[189], stage099[254]}
   );
   gpc606_5 gpc606_5_5761(
      {stage099[186], stage099[187], stage099[188], stage099[189], stage099[190], stage099[191]},
      {stage101[152], stage101[153], stage101[154], stage101[155], stage101[156], stage101[157]},
      {stage103[196], stage102[205], stage101[197], stage100[190], stage099[255]}
   );
   gpc606_5 gpc606_5_5762(
      {stage099[192], stage099[193], stage099[194], stage099[195], stage099[196], stage099[197]},
      {stage101[158], stage101[159], stage101[160], stage101[161], stage101[162], stage101[163]},
      {stage103[197], stage102[206], stage101[198], stage100[191], stage099[256]}
   );
   gpc606_5 gpc606_5_5763(
      {stage099[198], stage099[199], stage099[200], stage099[201], stage099[202], stage099[203]},
      {stage101[164], stage101[165], stage101[166], stage101[167], stage101[168], stage101[169]},
      {stage103[198], stage102[207], stage101[199], stage100[192], stage099[257]}
   );
   gpc1_1 gpc1_1_5764(
      {stage100[134]},
      {stage100[193]}
   );
   gpc1_1 gpc1_1_5765(
      {stage100[135]},
      {stage100[194]}
   );
   gpc606_5 gpc606_5_5766(
      {stage100[136], stage100[137], stage100[138], stage100[139], stage100[140], stage100[141]},
      {stage102[128], stage102[129], stage102[130], stage102[131], stage102[132], stage102[133]},
      {stage104[211], stage103[199], stage102[208], stage101[200], stage100[195]}
   );
   gpc606_5 gpc606_5_5767(
      {stage100[142], stage100[143], stage100[144], stage100[145], stage100[146], stage100[147]},
      {stage102[134], stage102[135], stage102[136], stage102[137], stage102[138], stage102[139]},
      {stage104[212], stage103[200], stage102[209], stage101[201], stage100[196]}
   );
   gpc606_5 gpc606_5_5768(
      {stage100[148], stage100[149], stage100[150], stage100[151], stage100[152], stage100[153]},
      {stage102[140], stage102[141], stage102[142], stage102[143], stage102[144], stage102[145]},
      {stage104[213], stage103[201], stage102[210], stage101[202], stage100[197]}
   );
   gpc606_5 gpc606_5_5769(
      {stage100[154], stage100[155], stage100[156], stage100[157], stage100[158], stage100[159]},
      {stage102[146], stage102[147], stage102[148], stage102[149], stage102[150], stage102[151]},
      {stage104[214], stage103[202], stage102[211], stage101[203], stage100[198]}
   );
   gpc606_5 gpc606_5_5770(
      {stage100[160], stage100[161], stage100[162], stage100[163], stage100[164], stage100[165]},
      {stage102[152], stage102[153], stage102[154], stage102[155], stage102[156], stage102[157]},
      {stage104[215], stage103[203], stage102[212], stage101[204], stage100[199]}
   );
   gpc606_5 gpc606_5_5771(
      {stage100[166], stage100[167], stage100[168], stage100[169], stage100[170], stage100[171]},
      {stage102[158], stage102[159], stage102[160], stage102[161], stage102[162], stage102[163]},
      {stage104[216], stage103[204], stage102[213], stage101[205], stage100[200]}
   );
   gpc606_5 gpc606_5_5772(
      {stage100[172], stage100[173], stage100[174], stage100[175], stage100[176], stage100[177]},
      {stage102[164], stage102[165], stage102[166], stage102[167], stage102[168], stage102[169]},
      {stage104[217], stage103[205], stage102[214], stage101[206], stage100[201]}
   );
   gpc1_1 gpc1_1_5773(
      {stage101[170]},
      {stage101[207]}
   );
   gpc1_1 gpc1_1_5774(
      {stage101[171]},
      {stage101[208]}
   );
   gpc1_1 gpc1_1_5775(
      {stage101[172]},
      {stage101[209]}
   );
   gpc1_1 gpc1_1_5776(
      {stage101[173]},
      {stage101[210]}
   );
   gpc1_1 gpc1_1_5777(
      {stage101[174]},
      {stage101[211]}
   );
   gpc1_1 gpc1_1_5778(
      {stage101[175]},
      {stage101[212]}
   );
   gpc1_1 gpc1_1_5779(
      {stage101[176]},
      {stage101[213]}
   );
   gpc1_1 gpc1_1_5780(
      {stage101[177]},
      {stage101[214]}
   );
   gpc1_1 gpc1_1_5781(
      {stage101[178]},
      {stage101[215]}
   );
   gpc1_1 gpc1_1_5782(
      {stage101[179]},
      {stage101[216]}
   );
   gpc1_1 gpc1_1_5783(
      {stage101[180]},
      {stage101[217]}
   );
   gpc1_1 gpc1_1_5784(
      {stage101[181]},
      {stage101[218]}
   );
   gpc1_1 gpc1_1_5785(
      {stage101[182]},
      {stage101[219]}
   );
   gpc1_1 gpc1_1_5786(
      {stage101[183]},
      {stage101[220]}
   );
   gpc1_1 gpc1_1_5787(
      {stage101[184]},
      {stage101[221]}
   );
   gpc1_1 gpc1_1_5788(
      {stage101[185]},
      {stage101[222]}
   );
   gpc1_1 gpc1_1_5789(
      {stage101[186]},
      {stage101[223]}
   );
   gpc1_1 gpc1_1_5790(
      {stage101[187]},
      {stage101[224]}
   );
   gpc1_1 gpc1_1_5791(
      {stage101[188]},
      {stage101[225]}
   );
   gpc1_1 gpc1_1_5792(
      {stage101[189]},
      {stage101[226]}
   );
   gpc1_1 gpc1_1_5793(
      {stage101[190]},
      {stage101[227]}
   );
   gpc1_1 gpc1_1_5794(
      {stage101[191]},
      {stage101[228]}
   );
   gpc615_5 gpc615_5_5795(
      {stage102[170], stage102[171], stage102[172], stage102[173], stage102[174]},
      {stage103[128]},
      {stage104[128], stage104[129], stage104[130], stage104[131], stage104[132], stage104[133]},
      {stage106[197], stage105[183], stage104[218], stage103[206], stage102[215]}
   );
   gpc615_5 gpc615_5_5796(
      {stage102[175], stage102[176], stage102[177], stage102[178], stage102[179]},
      {stage103[129]},
      {stage104[134], stage104[135], stage104[136], stage104[137], stage104[138], stage104[139]},
      {stage106[198], stage105[184], stage104[219], stage103[207], stage102[216]}
   );
   gpc615_5 gpc615_5_5797(
      {stage102[180], stage102[181], stage102[182], stage102[183], stage102[184]},
      {stage103[130]},
      {stage104[140], stage104[141], stage104[142], stage104[143], stage104[144], stage104[145]},
      {stage106[199], stage105[185], stage104[220], stage103[208], stage102[217]}
   );
   gpc615_5 gpc615_5_5798(
      {stage102[185], stage102[186], stage102[187], stage102[188], stage102[189]},
      {stage103[131]},
      {stage104[146], stage104[147], stage104[148], stage104[149], stage104[150], stage104[151]},
      {stage106[200], stage105[186], stage104[221], stage103[209], stage102[218]}
   );
   gpc615_5 gpc615_5_5799(
      {stage102[190], stage102[191], stage102[192], stage102[193], stage102[194]},
      {stage103[132]},
      {stage104[152], stage104[153], stage104[154], stage104[155], stage104[156], stage104[157]},
      {stage106[201], stage105[187], stage104[222], stage103[210], stage102[219]}
   );
   gpc615_5 gpc615_5_5800(
      {stage102[195], stage102[196], stage102[197], stage102[198], stage102[199]},
      {stage103[133]},
      {stage104[158], stage104[159], stage104[160], stage104[161], stage104[162], stage104[163]},
      {stage106[202], stage105[188], stage104[223], stage103[211], stage102[220]}
   );
   gpc1_1 gpc1_1_5801(
      {stage103[134]},
      {stage103[212]}
   );
   gpc1_1 gpc1_1_5802(
      {stage103[135]},
      {stage103[213]}
   );
   gpc1_1 gpc1_1_5803(
      {stage103[136]},
      {stage103[214]}
   );
   gpc1_1 gpc1_1_5804(
      {stage103[137]},
      {stage103[215]}
   );
   gpc606_5 gpc606_5_5805(
      {stage103[138], stage103[139], stage103[140], stage103[141], stage103[142], stage103[143]},
      {stage105[128], stage105[129], stage105[130], stage105[131], stage105[132], stage105[133]},
      {stage107[187], stage106[203], stage105[189], stage104[224], stage103[216]}
   );
   gpc606_5 gpc606_5_5806(
      {stage103[144], stage103[145], stage103[146], stage103[147], stage103[148], stage103[149]},
      {stage105[134], stage105[135], stage105[136], stage105[137], stage105[138], stage105[139]},
      {stage107[188], stage106[204], stage105[190], stage104[225], stage103[217]}
   );
   gpc606_5 gpc606_5_5807(
      {stage103[150], stage103[151], stage103[152], stage103[153], stage103[154], stage103[155]},
      {stage105[140], stage105[141], stage105[142], stage105[143], stage105[144], stage105[145]},
      {stage107[189], stage106[205], stage105[191], stage104[226], stage103[218]}
   );
   gpc606_5 gpc606_5_5808(
      {stage103[156], stage103[157], stage103[158], stage103[159], stage103[160], stage103[161]},
      {stage105[146], stage105[147], stage105[148], stage105[149], stage105[150], stage105[151]},
      {stage107[190], stage106[206], stage105[192], stage104[227], stage103[219]}
   );
   gpc606_5 gpc606_5_5809(
      {stage103[162], stage103[163], stage103[164], stage103[165], stage103[166], stage103[167]},
      {stage105[152], stage105[153], stage105[154], stage105[155], stage105[156], stage105[157]},
      {stage107[191], stage106[207], stage105[193], stage104[228], stage103[220]}
   );
   gpc606_5 gpc606_5_5810(
      {stage103[168], stage103[169], stage103[170], stage103[171], stage103[172], stage103[173]},
      {stage105[158], stage105[159], stage105[160], stage105[161], stage105[162], stage105[163]},
      {stage107[192], stage106[208], stage105[194], stage104[229], stage103[221]}
   );
   gpc606_5 gpc606_5_5811(
      {stage103[174], stage103[175], stage103[176], stage103[177], stage103[178], stage103[179]},
      {stage105[164], stage105[165], stage105[166], stage105[167], stage105[168], stage105[169]},
      {stage107[193], stage106[209], stage105[195], stage104[230], stage103[222]}
   );
   gpc606_5 gpc606_5_5812(
      {stage103[180], stage103[181], stage103[182], stage103[183], stage103[184], stage103[185]},
      {stage105[170], stage105[171], stage105[172], stage105[173], stage105[174], stage105[175]},
      {stage107[194], stage106[210], stage105[196], stage104[231], stage103[223]}
   );
   gpc606_5 gpc606_5_5813(
      {stage103[186], stage103[187], stage103[188], stage103[189], stage103[190], stage103[191]},
      {stage105[176], stage105[177], stage105[178], stage105[179], stage105[180], stage105[181]},
      {stage107[195], stage106[211], stage105[197], stage104[232], stage103[224]}
   );
   gpc1_1 gpc1_1_5814(
      {stage104[164]},
      {stage104[233]}
   );
   gpc1_1 gpc1_1_5815(
      {stage104[165]},
      {stage104[234]}
   );
   gpc1_1 gpc1_1_5816(
      {stage104[166]},
      {stage104[235]}
   );
   gpc1_1 gpc1_1_5817(
      {stage104[167]},
      {stage104[236]}
   );
   gpc1_1 gpc1_1_5818(
      {stage104[168]},
      {stage104[237]}
   );
   gpc606_5 gpc606_5_5819(
      {stage104[169], stage104[170], stage104[171], stage104[172], stage104[173], stage104[174]},
      {stage106[128], stage106[129], stage106[130], stage106[131], stage106[132], stage106[133]},
      {stage108[180], stage107[196], stage106[212], stage105[198], stage104[238]}
   );
   gpc606_5 gpc606_5_5820(
      {stage104[175], stage104[176], stage104[177], stage104[178], stage104[179], stage104[180]},
      {stage106[134], stage106[135], stage106[136], stage106[137], stage106[138], stage106[139]},
      {stage108[181], stage107[197], stage106[213], stage105[199], stage104[239]}
   );
   gpc606_5 gpc606_5_5821(
      {stage104[181], stage104[182], stage104[183], stage104[184], stage104[185], stage104[186]},
      {stage106[140], stage106[141], stage106[142], stage106[143], stage106[144], stage106[145]},
      {stage108[182], stage107[198], stage106[214], stage105[200], stage104[240]}
   );
   gpc606_5 gpc606_5_5822(
      {stage104[187], stage104[188], stage104[189], stage104[190], stage104[191], stage104[192]},
      {stage106[146], stage106[147], stage106[148], stage106[149], stage106[150], stage106[151]},
      {stage108[183], stage107[199], stage106[215], stage105[201], stage104[241]}
   );
   gpc606_5 gpc606_5_5823(
      {stage104[193], stage104[194], stage104[195], stage104[196], stage104[197], stage104[198]},
      {stage106[152], stage106[153], stage106[154], stage106[155], stage106[156], stage106[157]},
      {stage108[184], stage107[200], stage106[216], stage105[202], stage104[242]}
   );
   gpc606_5 gpc606_5_5824(
      {stage104[199], stage104[200], stage104[201], stage104[202], stage104[203], stage104[204]},
      {stage106[158], stage106[159], stage106[160], stage106[161], stage106[162], stage106[163]},
      {stage108[185], stage107[201], stage106[217], stage105[203], stage104[243]}
   );
   gpc606_5 gpc606_5_5825(
      {stage104[205], stage104[206], stage104[207], stage104[208], stage104[209], stage104[210]},
      {stage106[164], stage106[165], stage106[166], stage106[167], stage106[168], stage106[169]},
      {stage108[186], stage107[202], stage106[218], stage105[204], stage104[244]}
   );
   gpc1_1 gpc1_1_5826(
      {stage105[182]},
      {stage105[205]}
   );
   gpc1_1 gpc1_1_5827(
      {stage106[170]},
      {stage106[219]}
   );
   gpc1_1 gpc1_1_5828(
      {stage106[171]},
      {stage106[220]}
   );
   gpc1_1 gpc1_1_5829(
      {stage106[172]},
      {stage106[221]}
   );
   gpc1_1 gpc1_1_5830(
      {stage106[173]},
      {stage106[222]}
   );
   gpc1_1 gpc1_1_5831(
      {stage106[174]},
      {stage106[223]}
   );
   gpc1_1 gpc1_1_5832(
      {stage106[175]},
      {stage106[224]}
   );
   gpc606_5 gpc606_5_5833(
      {stage106[176], stage106[177], stage106[178], stage106[179], stage106[180], stage106[181]},
      {stage108[128], stage108[129], stage108[130], stage108[131], stage108[132], stage108[133]},
      {stage110[199], stage109[183], stage108[187], stage107[203], stage106[225]}
   );
   gpc615_5 gpc615_5_5834(
      {stage106[182], stage106[183], stage106[184], stage106[185], stage106[186]},
      {stage107[128]},
      {stage108[134], stage108[135], stage108[136], stage108[137], stage108[138], stage108[139]},
      {stage110[200], stage109[184], stage108[188], stage107[204], stage106[226]}
   );
   gpc615_5 gpc615_5_5835(
      {stage106[187], stage106[188], stage106[189], stage106[190], stage106[191]},
      {stage107[129]},
      {stage108[140], stage108[141], stage108[142], stage108[143], stage108[144], stage108[145]},
      {stage110[201], stage109[185], stage108[189], stage107[205], stage106[227]}
   );
   gpc615_5 gpc615_5_5836(
      {stage106[192], stage106[193], stage106[194], stage106[195], stage106[196]},
      {stage107[130]},
      {stage108[146], stage108[147], stage108[148], stage108[149], stage108[150], stage108[151]},
      {stage110[202], stage109[186], stage108[190], stage107[206], stage106[228]}
   );
   gpc1_1 gpc1_1_5837(
      {stage107[131]},
      {stage107[207]}
   );
   gpc1_1 gpc1_1_5838(
      {stage107[132]},
      {stage107[208]}
   );
   gpc1_1 gpc1_1_5839(
      {stage107[133]},
      {stage107[209]}
   );
   gpc1_1 gpc1_1_5840(
      {stage107[134]},
      {stage107[210]}
   );
   gpc1_1 gpc1_1_5841(
      {stage107[135]},
      {stage107[211]}
   );
   gpc1_1 gpc1_1_5842(
      {stage107[136]},
      {stage107[212]}
   );
   gpc1_1 gpc1_1_5843(
      {stage107[137]},
      {stage107[213]}
   );
   gpc1_1 gpc1_1_5844(
      {stage107[138]},
      {stage107[214]}
   );
   gpc1_1 gpc1_1_5845(
      {stage107[139]},
      {stage107[215]}
   );
   gpc1_1 gpc1_1_5846(
      {stage107[140]},
      {stage107[216]}
   );
   gpc1_1 gpc1_1_5847(
      {stage107[141]},
      {stage107[217]}
   );
   gpc1_1 gpc1_1_5848(
      {stage107[142]},
      {stage107[218]}
   );
   gpc1_1 gpc1_1_5849(
      {stage107[143]},
      {stage107[219]}
   );
   gpc1_1 gpc1_1_5850(
      {stage107[144]},
      {stage107[220]}
   );
   gpc1_1 gpc1_1_5851(
      {stage107[145]},
      {stage107[221]}
   );
   gpc7_3 gpc7_3_5852(
      {stage107[146], stage107[147], stage107[148], stage107[149], stage107[150], stage107[151], stage107[152]},
      {stage109[187], stage108[191], stage107[222]}
   );
   gpc7_3 gpc7_3_5853(
      {stage107[153], stage107[154], stage107[155], stage107[156], stage107[157], stage107[158], stage107[159]},
      {stage109[188], stage108[192], stage107[223]}
   );
   gpc7_3 gpc7_3_5854(
      {stage107[160], stage107[161], stage107[162], stage107[163], stage107[164], stage107[165], stage107[166]},
      {stage109[189], stage108[193], stage107[224]}
   );
   gpc7_3 gpc7_3_5855(
      {stage107[167], stage107[168], stage107[169], stage107[170], stage107[171], stage107[172], stage107[173]},
      {stage109[190], stage108[194], stage107[225]}
   );
   gpc7_3 gpc7_3_5856(
      {stage107[174], stage107[175], stage107[176], stage107[177], stage107[178], stage107[179], stage107[180]},
      {stage109[191], stage108[195], stage107[226]}
   );
   gpc606_5 gpc606_5_5857(
      {stage107[181], stage107[182], stage107[183], stage107[184], stage107[185], stage107[186]},
      {stage109[128], stage109[129], stage109[130], stage109[131], stage109[132], stage109[133]},
      {stage111[215], stage110[203], stage109[192], stage108[196], stage107[227]}
   );
   gpc1_1 gpc1_1_5858(
      {stage108[152]},
      {stage108[197]}
   );
   gpc1_1 gpc1_1_5859(
      {stage108[153]},
      {stage108[198]}
   );
   gpc1_1 gpc1_1_5860(
      {stage108[154]},
      {stage108[199]}
   );
   gpc1_1 gpc1_1_5861(
      {stage108[155]},
      {stage108[200]}
   );
   gpc1_1 gpc1_1_5862(
      {stage108[156]},
      {stage108[201]}
   );
   gpc1_1 gpc1_1_5863(
      {stage108[157]},
      {stage108[202]}
   );
   gpc1_1 gpc1_1_5864(
      {stage108[158]},
      {stage108[203]}
   );
   gpc1_1 gpc1_1_5865(
      {stage108[159]},
      {stage108[204]}
   );
   gpc1_1 gpc1_1_5866(
      {stage108[160]},
      {stage108[205]}
   );
   gpc1_1 gpc1_1_5867(
      {stage108[161]},
      {stage108[206]}
   );
   gpc1_1 gpc1_1_5868(
      {stage108[162]},
      {stage108[207]}
   );
   gpc1_1 gpc1_1_5869(
      {stage108[163]},
      {stage108[208]}
   );
   gpc1_1 gpc1_1_5870(
      {stage108[164]},
      {stage108[209]}
   );
   gpc1_1 gpc1_1_5871(
      {stage108[165]},
      {stage108[210]}
   );
   gpc1_1 gpc1_1_5872(
      {stage108[166]},
      {stage108[211]}
   );
   gpc1_1 gpc1_1_5873(
      {stage108[167]},
      {stage108[212]}
   );
   gpc1_1 gpc1_1_5874(
      {stage108[168]},
      {stage108[213]}
   );
   gpc1_1 gpc1_1_5875(
      {stage108[169]},
      {stage108[214]}
   );
   gpc1_1 gpc1_1_5876(
      {stage108[170]},
      {stage108[215]}
   );
   gpc1_1 gpc1_1_5877(
      {stage108[171]},
      {stage108[216]}
   );
   gpc1_1 gpc1_1_5878(
      {stage108[172]},
      {stage108[217]}
   );
   gpc1_1 gpc1_1_5879(
      {stage108[173]},
      {stage108[218]}
   );
   gpc1_1 gpc1_1_5880(
      {stage108[174]},
      {stage108[219]}
   );
   gpc1_1 gpc1_1_5881(
      {stage108[175]},
      {stage108[220]}
   );
   gpc1_1 gpc1_1_5882(
      {stage108[176]},
      {stage108[221]}
   );
   gpc1_1 gpc1_1_5883(
      {stage108[177]},
      {stage108[222]}
   );
   gpc1_1 gpc1_1_5884(
      {stage108[178]},
      {stage108[223]}
   );
   gpc1_1 gpc1_1_5885(
      {stage108[179]},
      {stage108[224]}
   );
   gpc1_1 gpc1_1_5886(
      {stage109[134]},
      {stage109[193]}
   );
   gpc1_1 gpc1_1_5887(
      {stage109[135]},
      {stage109[194]}
   );
   gpc1_1 gpc1_1_5888(
      {stage109[136]},
      {stage109[195]}
   );
   gpc1_1 gpc1_1_5889(
      {stage109[137]},
      {stage109[196]}
   );
   gpc1_1 gpc1_1_5890(
      {stage109[138]},
      {stage109[197]}
   );
   gpc1_1 gpc1_1_5891(
      {stage109[139]},
      {stage109[198]}
   );
   gpc1_1 gpc1_1_5892(
      {stage109[140]},
      {stage109[199]}
   );
   gpc1_1 gpc1_1_5893(
      {stage109[141]},
      {stage109[200]}
   );
   gpc606_5 gpc606_5_5894(
      {stage109[142], stage109[143], stage109[144], stage109[145], stage109[146], stage109[147]},
      {stage111[128], stage111[129], stage111[130], stage111[131], stage111[132], stage111[133]},
      {stage113[183], stage112[192], stage111[216], stage110[204], stage109[201]}
   );
   gpc615_5 gpc615_5_5895(
      {stage109[148], stage109[149], stage109[150], stage109[151], stage109[152]},
      {stage110[128]},
      {stage111[134], stage111[135], stage111[136], stage111[137], stage111[138], stage111[139]},
      {stage113[184], stage112[193], stage111[217], stage110[205], stage109[202]}
   );
   gpc615_5 gpc615_5_5896(
      {stage109[153], stage109[154], stage109[155], stage109[156], stage109[157]},
      {stage110[129]},
      {stage111[140], stage111[141], stage111[142], stage111[143], stage111[144], stage111[145]},
      {stage113[185], stage112[194], stage111[218], stage110[206], stage109[203]}
   );
   gpc615_5 gpc615_5_5897(
      {stage109[158], stage109[159], stage109[160], stage109[161], stage109[162]},
      {stage110[130]},
      {stage111[146], stage111[147], stage111[148], stage111[149], stage111[150], stage111[151]},
      {stage113[186], stage112[195], stage111[219], stage110[207], stage109[204]}
   );
   gpc615_5 gpc615_5_5898(
      {stage109[163], stage109[164], stage109[165], stage109[166], stage109[167]},
      {stage110[131]},
      {stage111[152], stage111[153], stage111[154], stage111[155], stage111[156], stage111[157]},
      {stage113[187], stage112[196], stage111[220], stage110[208], stage109[205]}
   );
   gpc615_5 gpc615_5_5899(
      {stage109[168], stage109[169], stage109[170], stage109[171], stage109[172]},
      {stage110[132]},
      {stage111[158], stage111[159], stage111[160], stage111[161], stage111[162], stage111[163]},
      {stage113[188], stage112[197], stage111[221], stage110[209], stage109[206]}
   );
   gpc615_5 gpc615_5_5900(
      {stage109[173], stage109[174], stage109[175], stage109[176], stage109[177]},
      {stage110[133]},
      {stage111[164], stage111[165], stage111[166], stage111[167], stage111[168], stage111[169]},
      {stage113[189], stage112[198], stage111[222], stage110[210], stage109[207]}
   );
   gpc615_5 gpc615_5_5901(
      {stage109[178], stage109[179], stage109[180], stage109[181], stage109[182]},
      {stage110[134]},
      {stage111[170], stage111[171], stage111[172], stage111[173], stage111[174], stage111[175]},
      {stage113[190], stage112[199], stage111[223], stage110[211], stage109[208]}
   );
   gpc1_1 gpc1_1_5902(
      {stage110[135]},
      {stage110[212]}
   );
   gpc1_1 gpc1_1_5903(
      {stage110[136]},
      {stage110[213]}
   );
   gpc1_1 gpc1_1_5904(
      {stage110[137]},
      {stage110[214]}
   );
   gpc1_1 gpc1_1_5905(
      {stage110[138]},
      {stage110[215]}
   );
   gpc1_1 gpc1_1_5906(
      {stage110[139]},
      {stage110[216]}
   );
   gpc1_1 gpc1_1_5907(
      {stage110[140]},
      {stage110[217]}
   );
   gpc1_1 gpc1_1_5908(
      {stage110[141]},
      {stage110[218]}
   );
   gpc1_1 gpc1_1_5909(
      {stage110[142]},
      {stage110[219]}
   );
   gpc1_1 gpc1_1_5910(
      {stage110[143]},
      {stage110[220]}
   );
   gpc1_1 gpc1_1_5911(
      {stage110[144]},
      {stage110[221]}
   );
   gpc1_1 gpc1_1_5912(
      {stage110[145]},
      {stage110[222]}
   );
   gpc1_1 gpc1_1_5913(
      {stage110[146]},
      {stage110[223]}
   );
   gpc1_1 gpc1_1_5914(
      {stage110[147]},
      {stage110[224]}
   );
   gpc1_1 gpc1_1_5915(
      {stage110[148]},
      {stage110[225]}
   );
   gpc615_5 gpc615_5_5916(
      {stage110[149], stage110[150], stage110[151], stage110[152], stage110[153]},
      {stage111[176]},
      {stage112[128], stage112[129], stage112[130], stage112[131], stage112[132], stage112[133]},
      {stage114[183], stage113[191], stage112[200], stage111[224], stage110[226]}
   );
   gpc615_5 gpc615_5_5917(
      {stage110[154], stage110[155], stage110[156], stage110[157], stage110[158]},
      {stage111[177]},
      {stage112[134], stage112[135], stage112[136], stage112[137], stage112[138], stage112[139]},
      {stage114[184], stage113[192], stage112[201], stage111[225], stage110[227]}
   );
   gpc615_5 gpc615_5_5918(
      {stage110[159], stage110[160], stage110[161], stage110[162], stage110[163]},
      {stage111[178]},
      {stage112[140], stage112[141], stage112[142], stage112[143], stage112[144], stage112[145]},
      {stage114[185], stage113[193], stage112[202], stage111[226], stage110[228]}
   );
   gpc615_5 gpc615_5_5919(
      {stage110[164], stage110[165], stage110[166], stage110[167], stage110[168]},
      {stage111[179]},
      {stage112[146], stage112[147], stage112[148], stage112[149], stage112[150], stage112[151]},
      {stage114[186], stage113[194], stage112[203], stage111[227], stage110[229]}
   );
   gpc615_5 gpc615_5_5920(
      {stage110[169], stage110[170], stage110[171], stage110[172], stage110[173]},
      {stage111[180]},
      {stage112[152], stage112[153], stage112[154], stage112[155], stage112[156], stage112[157]},
      {stage114[187], stage113[195], stage112[204], stage111[228], stage110[230]}
   );
   gpc615_5 gpc615_5_5921(
      {stage110[174], stage110[175], stage110[176], stage110[177], stage110[178]},
      {stage111[181]},
      {stage112[158], stage112[159], stage112[160], stage112[161], stage112[162], stage112[163]},
      {stage114[188], stage113[196], stage112[205], stage111[229], stage110[231]}
   );
   gpc615_5 gpc615_5_5922(
      {stage110[179], stage110[180], stage110[181], stage110[182], stage110[183]},
      {stage111[182]},
      {stage112[164], stage112[165], stage112[166], stage112[167], stage112[168], stage112[169]},
      {stage114[189], stage113[197], stage112[206], stage111[230], stage110[232]}
   );
   gpc615_5 gpc615_5_5923(
      {stage110[184], stage110[185], stage110[186], stage110[187], stage110[188]},
      {stage111[183]},
      {stage112[170], stage112[171], stage112[172], stage112[173], stage112[174], stage112[175]},
      {stage114[190], stage113[198], stage112[207], stage111[231], stage110[233]}
   );
   gpc615_5 gpc615_5_5924(
      {stage110[189], stage110[190], stage110[191], stage110[192], stage110[193]},
      {stage111[184]},
      {stage112[176], stage112[177], stage112[178], stage112[179], stage112[180], stage112[181]},
      {stage114[191], stage113[199], stage112[208], stage111[232], stage110[234]}
   );
   gpc615_5 gpc615_5_5925(
      {stage110[194], stage110[195], stage110[196], stage110[197], stage110[198]},
      {stage111[185]},
      {stage112[182], stage112[183], stage112[184], stage112[185], stage112[186], stage112[187]},
      {stage114[192], stage113[200], stage112[209], stage111[233], stage110[235]}
   );
   gpc1_1 gpc1_1_5926(
      {stage111[186]},
      {stage111[234]}
   );
   gpc1_1 gpc1_1_5927(
      {stage111[187]},
      {stage111[235]}
   );
   gpc1_1 gpc1_1_5928(
      {stage111[188]},
      {stage111[236]}
   );
   gpc615_5 gpc615_5_5929(
      {stage111[189], stage111[190], stage111[191], stage111[192], stage111[193]},
      {stage112[188]},
      {stage113[128], stage113[129], stage113[130], stage113[131], stage113[132], stage113[133]},
      {stage115[196], stage114[193], stage113[201], stage112[210], stage111[237]}
   );
   gpc615_5 gpc615_5_5930(
      {stage111[194], stage111[195], stage111[196], stage111[197], stage111[198]},
      {stage112[189]},
      {stage113[134], stage113[135], stage113[136], stage113[137], stage113[138], stage113[139]},
      {stage115[197], stage114[194], stage113[202], stage112[211], stage111[238]}
   );
   gpc615_5 gpc615_5_5931(
      {stage111[199], stage111[200], stage111[201], stage111[202], stage111[203]},
      {stage112[190]},
      {stage113[140], stage113[141], stage113[142], stage113[143], stage113[144], stage113[145]},
      {stage115[198], stage114[195], stage113[203], stage112[212], stage111[239]}
   );
   gpc615_5 gpc615_5_5932(
      {stage111[204], stage111[205], stage111[206], stage111[207], stage111[208]},
      {stage112[191]},
      {stage113[146], stage113[147], stage113[148], stage113[149], stage113[150], stage113[151]},
      {stage115[199], stage114[196], stage113[204], stage112[213], stage111[240]}
   );
   gpc1406_5 gpc1406_5_5933(
      {stage111[209], stage111[210], stage111[211], stage111[212], stage111[213], stage111[214]},
      {stage113[152], stage113[153], stage113[154], stage113[155]},
      {stage114[128]},
      {stage115[200], stage114[197], stage113[205], stage112[214], stage111[241]}
   );
   gpc1_1 gpc1_1_5934(
      {stage113[156]},
      {stage113[206]}
   );
   gpc1_1 gpc1_1_5935(
      {stage113[157]},
      {stage113[207]}
   );
   gpc1_1 gpc1_1_5936(
      {stage113[158]},
      {stage113[208]}
   );
   gpc606_5 gpc606_5_5937(
      {stage113[159], stage113[160], stage113[161], stage113[162], stage113[163], stage113[164]},
      {stage115[128], stage115[129], stage115[130], stage115[131], stage115[132], stage115[133]},
      {stage117[196], stage116[187], stage115[201], stage114[198], stage113[209]}
   );
   gpc606_5 gpc606_5_5938(
      {stage113[165], stage113[166], stage113[167], stage113[168], stage113[169], stage113[170]},
      {stage115[134], stage115[135], stage115[136], stage115[137], stage115[138], stage115[139]},
      {stage117[197], stage116[188], stage115[202], stage114[199], stage113[210]}
   );
   gpc606_5 gpc606_5_5939(
      {stage113[171], stage113[172], stage113[173], stage113[174], stage113[175], stage113[176]},
      {stage115[140], stage115[141], stage115[142], stage115[143], stage115[144], stage115[145]},
      {stage117[198], stage116[189], stage115[203], stage114[200], stage113[211]}
   );
   gpc606_5 gpc606_5_5940(
      {stage113[177], stage113[178], stage113[179], stage113[180], stage113[181], stage113[182]},
      {stage115[146], stage115[147], stage115[148], stage115[149], stage115[150], stage115[151]},
      {stage117[199], stage116[190], stage115[204], stage114[201], stage113[212]}
   );
   gpc1_1 gpc1_1_5941(
      {stage114[129]},
      {stage114[202]}
   );
   gpc1_1 gpc1_1_5942(
      {stage114[130]},
      {stage114[203]}
   );
   gpc1_1 gpc1_1_5943(
      {stage114[131]},
      {stage114[204]}
   );
   gpc1_1 gpc1_1_5944(
      {stage114[132]},
      {stage114[205]}
   );
   gpc1_1 gpc1_1_5945(
      {stage114[133]},
      {stage114[206]}
   );
   gpc1_1 gpc1_1_5946(
      {stage114[134]},
      {stage114[207]}
   );
   gpc606_5 gpc606_5_5947(
      {stage114[135], stage114[136], stage114[137], stage114[138], stage114[139], stage114[140]},
      {stage116[128], stage116[129], stage116[130], stage116[131], stage116[132], stage116[133]},
      {stage118[183], stage117[200], stage116[191], stage115[205], stage114[208]}
   );
   gpc606_5 gpc606_5_5948(
      {stage114[141], stage114[142], stage114[143], stage114[144], stage114[145], stage114[146]},
      {stage116[134], stage116[135], stage116[136], stage116[137], stage116[138], stage116[139]},
      {stage118[184], stage117[201], stage116[192], stage115[206], stage114[209]}
   );
   gpc606_5 gpc606_5_5949(
      {stage114[147], stage114[148], stage114[149], stage114[150], stage114[151], stage114[152]},
      {stage116[140], stage116[141], stage116[142], stage116[143], stage116[144], stage116[145]},
      {stage118[185], stage117[202], stage116[193], stage115[207], stage114[210]}
   );
   gpc606_5 gpc606_5_5950(
      {stage114[153], stage114[154], stage114[155], stage114[156], stage114[157], stage114[158]},
      {stage116[146], stage116[147], stage116[148], stage116[149], stage116[150], stage116[151]},
      {stage118[186], stage117[203], stage116[194], stage115[208], stage114[211]}
   );
   gpc606_5 gpc606_5_5951(
      {stage114[159], stage114[160], stage114[161], stage114[162], stage114[163], stage114[164]},
      {stage116[152], stage116[153], stage116[154], stage116[155], stage116[156], stage116[157]},
      {stage118[187], stage117[204], stage116[195], stage115[209], stage114[212]}
   );
   gpc606_5 gpc606_5_5952(
      {stage114[165], stage114[166], stage114[167], stage114[168], stage114[169], stage114[170]},
      {stage116[158], stage116[159], stage116[160], stage116[161], stage116[162], stage116[163]},
      {stage118[188], stage117[205], stage116[196], stage115[210], stage114[213]}
   );
   gpc606_5 gpc606_5_5953(
      {stage114[171], stage114[172], stage114[173], stage114[174], stage114[175], stage114[176]},
      {stage116[164], stage116[165], stage116[166], stage116[167], stage116[168], stage116[169]},
      {stage118[189], stage117[206], stage116[197], stage115[211], stage114[214]}
   );
   gpc1406_5 gpc1406_5_5954(
      {stage114[177], stage114[178], stage114[179], stage114[180], stage114[181], stage114[182]},
      {stage116[170], stage116[171], stage116[172], stage116[173]},
      {stage117[128]},
      {stage118[190], stage117[207], stage116[198], stage115[212], stage114[215]}
   );
   gpc1_1 gpc1_1_5955(
      {stage115[152]},
      {stage115[213]}
   );
   gpc1_1 gpc1_1_5956(
      {stage115[153]},
      {stage115[214]}
   );
   gpc1_1 gpc1_1_5957(
      {stage115[154]},
      {stage115[215]}
   );
   gpc1_1 gpc1_1_5958(
      {stage115[155]},
      {stage115[216]}
   );
   gpc1_1 gpc1_1_5959(
      {stage115[156]},
      {stage115[217]}
   );
   gpc1_1 gpc1_1_5960(
      {stage115[157]},
      {stage115[218]}
   );
   gpc1_1 gpc1_1_5961(
      {stage115[158]},
      {stage115[219]}
   );
   gpc1_1 gpc1_1_5962(
      {stage115[159]},
      {stage115[220]}
   );
   gpc1_1 gpc1_1_5963(
      {stage115[160]},
      {stage115[221]}
   );
   gpc1_1 gpc1_1_5964(
      {stage115[161]},
      {stage115[222]}
   );
   gpc1_1 gpc1_1_5965(
      {stage115[162]},
      {stage115[223]}
   );
   gpc1_1 gpc1_1_5966(
      {stage115[163]},
      {stage115[224]}
   );
   gpc1_1 gpc1_1_5967(
      {stage115[164]},
      {stage115[225]}
   );
   gpc1_1 gpc1_1_5968(
      {stage115[165]},
      {stage115[226]}
   );
   gpc1_1 gpc1_1_5969(
      {stage115[166]},
      {stage115[227]}
   );
   gpc1_1 gpc1_1_5970(
      {stage115[167]},
      {stage115[228]}
   );
   gpc1_1 gpc1_1_5971(
      {stage115[168]},
      {stage115[229]}
   );
   gpc1_1 gpc1_1_5972(
      {stage115[169]},
      {stage115[230]}
   );
   gpc1_1 gpc1_1_5973(
      {stage115[170]},
      {stage115[231]}
   );
   gpc1_1 gpc1_1_5974(
      {stage115[171]},
      {stage115[232]}
   );
   gpc606_5 gpc606_5_5975(
      {stage115[172], stage115[173], stage115[174], stage115[175], stage115[176], stage115[177]},
      {stage117[129], stage117[130], stage117[131], stage117[132], stage117[133], stage117[134]},
      {stage119[184], stage118[191], stage117[208], stage116[199], stage115[233]}
   );
   gpc606_5 gpc606_5_5976(
      {stage115[178], stage115[179], stage115[180], stage115[181], stage115[182], stage115[183]},
      {stage117[135], stage117[136], stage117[137], stage117[138], stage117[139], stage117[140]},
      {stage119[185], stage118[192], stage117[209], stage116[200], stage115[234]}
   );
   gpc606_5 gpc606_5_5977(
      {stage115[184], stage115[185], stage115[186], stage115[187], stage115[188], stage115[189]},
      {stage117[141], stage117[142], stage117[143], stage117[144], stage117[145], stage117[146]},
      {stage119[186], stage118[193], stage117[210], stage116[201], stage115[235]}
   );
   gpc606_5 gpc606_5_5978(
      {stage115[190], stage115[191], stage115[192], stage115[193], stage115[194], stage115[195]},
      {stage117[147], stage117[148], stage117[149], stage117[150], stage117[151], stage117[152]},
      {stage119[187], stage118[194], stage117[211], stage116[202], stage115[236]}
   );
   gpc1_1 gpc1_1_5979(
      {stage116[174]},
      {stage116[203]}
   );
   gpc1_1 gpc1_1_5980(
      {stage116[175]},
      {stage116[204]}
   );
   gpc1_1 gpc1_1_5981(
      {stage116[176]},
      {stage116[205]}
   );
   gpc1_1 gpc1_1_5982(
      {stage116[177]},
      {stage116[206]}
   );
   gpc1_1 gpc1_1_5983(
      {stage116[178]},
      {stage116[207]}
   );
   gpc1_1 gpc1_1_5984(
      {stage116[179]},
      {stage116[208]}
   );
   gpc1_1 gpc1_1_5985(
      {stage116[180]},
      {stage116[209]}
   );
   gpc1_1 gpc1_1_5986(
      {stage116[181]},
      {stage116[210]}
   );
   gpc1_1 gpc1_1_5987(
      {stage116[182]},
      {stage116[211]}
   );
   gpc1_1 gpc1_1_5988(
      {stage116[183]},
      {stage116[212]}
   );
   gpc623_5 gpc623_5_5989(
      {stage116[184], stage116[185], stage116[186]},
      {stage117[153], stage117[154]},
      {stage118[128], stage118[129], stage118[130], stage118[131], stage118[132], stage118[133]},
      {stage120[185], stage119[188], stage118[195], stage117[212], stage116[213]}
   );
   gpc1_1 gpc1_1_5990(
      {stage117[155]},
      {stage117[213]}
   );
   gpc1_1 gpc1_1_5991(
      {stage117[156]},
      {stage117[214]}
   );
   gpc1_1 gpc1_1_5992(
      {stage117[157]},
      {stage117[215]}
   );
   gpc606_5 gpc606_5_5993(
      {stage117[158], stage117[159], stage117[160], stage117[161], stage117[162], stage117[163]},
      {stage119[128], stage119[129], stage119[130], stage119[131], stage119[132], stage119[133]},
      {stage121[176], stage120[186], stage119[189], stage118[196], stage117[216]}
   );
   gpc606_5 gpc606_5_5994(
      {stage117[164], stage117[165], stage117[166], stage117[167], stage117[168], stage117[169]},
      {stage119[134], stage119[135], stage119[136], stage119[137], stage119[138], stage119[139]},
      {stage121[177], stage120[187], stage119[190], stage118[197], stage117[217]}
   );
   gpc606_5 gpc606_5_5995(
      {stage117[170], stage117[171], stage117[172], stage117[173], stage117[174], stage117[175]},
      {stage119[140], stage119[141], stage119[142], stage119[143], stage119[144], stage119[145]},
      {stage121[178], stage120[188], stage119[191], stage118[198], stage117[218]}
   );
   gpc615_5 gpc615_5_5996(
      {stage117[176], stage117[177], stage117[178], stage117[179], stage117[180]},
      {stage118[134]},
      {stage119[146], stage119[147], stage119[148], stage119[149], stage119[150], stage119[151]},
      {stage121[179], stage120[189], stage119[192], stage118[199], stage117[219]}
   );
   gpc615_5 gpc615_5_5997(
      {stage117[181], stage117[182], stage117[183], stage117[184], stage117[185]},
      {stage118[135]},
      {stage119[152], stage119[153], stage119[154], stage119[155], stage119[156], stage119[157]},
      {stage121[180], stage120[190], stage119[193], stage118[200], stage117[220]}
   );
   gpc615_5 gpc615_5_5998(
      {stage117[186], stage117[187], stage117[188], stage117[189], stage117[190]},
      {stage118[136]},
      {stage119[158], stage119[159], stage119[160], stage119[161], stage119[162], stage119[163]},
      {stage121[181], stage120[191], stage119[194], stage118[201], stage117[221]}
   );
   gpc615_5 gpc615_5_5999(
      {stage117[191], stage117[192], stage117[193], stage117[194], stage117[195]},
      {stage118[137]},
      {stage119[164], stage119[165], stage119[166], stage119[167], stage119[168], stage119[169]},
      {stage121[182], stage120[192], stage119[195], stage118[202], stage117[222]}
   );
   gpc1_1 gpc1_1_6000(
      {stage118[138]},
      {stage118[203]}
   );
   gpc1_1 gpc1_1_6001(
      {stage118[139]},
      {stage118[204]}
   );
   gpc1_1 gpc1_1_6002(
      {stage118[140]},
      {stage118[205]}
   );
   gpc1_1 gpc1_1_6003(
      {stage118[141]},
      {stage118[206]}
   );
   gpc1_1 gpc1_1_6004(
      {stage118[142]},
      {stage118[207]}
   );
   gpc1_1 gpc1_1_6005(
      {stage118[143]},
      {stage118[208]}
   );
   gpc1_1 gpc1_1_6006(
      {stage118[144]},
      {stage118[209]}
   );
   gpc1_1 gpc1_1_6007(
      {stage118[145]},
      {stage118[210]}
   );
   gpc1_1 gpc1_1_6008(
      {stage118[146]},
      {stage118[211]}
   );
   gpc1_1 gpc1_1_6009(
      {stage118[147]},
      {stage118[212]}
   );
   gpc1_1 gpc1_1_6010(
      {stage118[148]},
      {stage118[213]}
   );
   gpc1_1 gpc1_1_6011(
      {stage118[149]},
      {stage118[214]}
   );
   gpc1_1 gpc1_1_6012(
      {stage118[150]},
      {stage118[215]}
   );
   gpc1_1 gpc1_1_6013(
      {stage118[151]},
      {stage118[216]}
   );
   gpc1_1 gpc1_1_6014(
      {stage118[152]},
      {stage118[217]}
   );
   gpc615_5 gpc615_5_6015(
      {stage118[153], stage118[154], stage118[155], stage118[156], stage118[157]},
      {stage119[170]},
      {stage120[128], stage120[129], stage120[130], stage120[131], stage120[132], stage120[133]},
      {stage122[187], stage121[183], stage120[193], stage119[196], stage118[218]}
   );
   gpc615_5 gpc615_5_6016(
      {stage118[158], stage118[159], stage118[160], stage118[161], stage118[162]},
      {stage119[171]},
      {stage120[134], stage120[135], stage120[136], stage120[137], stage120[138], stage120[139]},
      {stage122[188], stage121[184], stage120[194], stage119[197], stage118[219]}
   );
   gpc615_5 gpc615_5_6017(
      {stage118[163], stage118[164], stage118[165], stage118[166], stage118[167]},
      {stage119[172]},
      {stage120[140], stage120[141], stage120[142], stage120[143], stage120[144], stage120[145]},
      {stage122[189], stage121[185], stage120[195], stage119[198], stage118[220]}
   );
   gpc615_5 gpc615_5_6018(
      {stage118[168], stage118[169], stage118[170], stage118[171], stage118[172]},
      {stage119[173]},
      {stage120[146], stage120[147], stage120[148], stage120[149], stage120[150], stage120[151]},
      {stage122[190], stage121[186], stage120[196], stage119[199], stage118[221]}
   );
   gpc615_5 gpc615_5_6019(
      {stage118[173], stage118[174], stage118[175], stage118[176], stage118[177]},
      {stage119[174]},
      {stage120[152], stage120[153], stage120[154], stage120[155], stage120[156], stage120[157]},
      {stage122[191], stage121[187], stage120[197], stage119[200], stage118[222]}
   );
   gpc615_5 gpc615_5_6020(
      {stage118[178], stage118[179], stage118[180], stage118[181], stage118[182]},
      {stage119[175]},
      {stage120[158], stage120[159], stage120[160], stage120[161], stage120[162], stage120[163]},
      {stage122[192], stage121[188], stage120[198], stage119[201], stage118[223]}
   );
   gpc1_1 gpc1_1_6021(
      {stage119[176]},
      {stage119[202]}
   );
   gpc1_1 gpc1_1_6022(
      {stage119[177]},
      {stage119[203]}
   );
   gpc1_1 gpc1_1_6023(
      {stage119[178]},
      {stage119[204]}
   );
   gpc1_1 gpc1_1_6024(
      {stage119[179]},
      {stage119[205]}
   );
   gpc1_1 gpc1_1_6025(
      {stage119[180]},
      {stage119[206]}
   );
   gpc1_1 gpc1_1_6026(
      {stage119[181]},
      {stage119[207]}
   );
   gpc1_1 gpc1_1_6027(
      {stage119[182]},
      {stage119[208]}
   );
   gpc1_1 gpc1_1_6028(
      {stage119[183]},
      {stage119[209]}
   );
   gpc1_1 gpc1_1_6029(
      {stage120[164]},
      {stage120[199]}
   );
   gpc1_1 gpc1_1_6030(
      {stage120[165]},
      {stage120[200]}
   );
   gpc1_1 gpc1_1_6031(
      {stage120[166]},
      {stage120[201]}
   );
   gpc1_1 gpc1_1_6032(
      {stage120[167]},
      {stage120[202]}
   );
   gpc1_1 gpc1_1_6033(
      {stage120[168]},
      {stage120[203]}
   );
   gpc1_1 gpc1_1_6034(
      {stage120[169]},
      {stage120[204]}
   );
   gpc1_1 gpc1_1_6035(
      {stage120[170]},
      {stage120[205]}
   );
   gpc1_1 gpc1_1_6036(
      {stage120[171]},
      {stage120[206]}
   );
   gpc1_1 gpc1_1_6037(
      {stage120[172]},
      {stage120[207]}
   );
   gpc1_1 gpc1_1_6038(
      {stage120[173]},
      {stage120[208]}
   );
   gpc1_1 gpc1_1_6039(
      {stage120[174]},
      {stage120[209]}
   );
   gpc1_1 gpc1_1_6040(
      {stage120[175]},
      {stage120[210]}
   );
   gpc1_1 gpc1_1_6041(
      {stage120[176]},
      {stage120[211]}
   );
   gpc1_1 gpc1_1_6042(
      {stage120[177]},
      {stage120[212]}
   );
   gpc1_1 gpc1_1_6043(
      {stage120[178]},
      {stage120[213]}
   );
   gpc1_1 gpc1_1_6044(
      {stage120[179]},
      {stage120[214]}
   );
   gpc1_1 gpc1_1_6045(
      {stage120[180]},
      {stage120[215]}
   );
   gpc1_1 gpc1_1_6046(
      {stage120[181]},
      {stage120[216]}
   );
   gpc1_1 gpc1_1_6047(
      {stage120[182]},
      {stage120[217]}
   );
   gpc1_1 gpc1_1_6048(
      {stage120[183]},
      {stage120[218]}
   );
   gpc1_1 gpc1_1_6049(
      {stage120[184]},
      {stage120[219]}
   );
   gpc1_1 gpc1_1_6050(
      {stage121[128]},
      {stage121[189]}
   );
   gpc1_1 gpc1_1_6051(
      {stage121[129]},
      {stage121[190]}
   );
   gpc1_1 gpc1_1_6052(
      {stage121[130]},
      {stage121[191]}
   );
   gpc1_1 gpc1_1_6053(
      {stage121[131]},
      {stage121[192]}
   );
   gpc1_1 gpc1_1_6054(
      {stage121[132]},
      {stage121[193]}
   );
   gpc1_1 gpc1_1_6055(
      {stage121[133]},
      {stage121[194]}
   );
   gpc1_1 gpc1_1_6056(
      {stage121[134]},
      {stage121[195]}
   );
   gpc623_5 gpc623_5_6057(
      {stage121[135], stage121[136], stage121[137]},
      {stage122[128], stage122[129]},
      {stage123[128], stage123[129], stage123[130], stage123[131], stage123[132], stage123[133]},
      {stage125[205], stage124[178], stage123[256], stage122[193], stage121[196]}
   );
   gpc623_5 gpc623_5_6058(
      {stage121[138], stage121[139], stage121[140]},
      {stage122[130], stage122[131]},
      {stage123[134], stage123[135], stage123[136], stage123[137], stage123[138], stage123[139]},
      {stage125[206], stage124[179], stage123[257], stage122[194], stage121[197]}
   );
   gpc615_5 gpc615_5_6059(
      {stage121[141], stage121[142], stage121[143], stage121[144], stage121[145]},
      {stage122[132]},
      {stage123[140], stage123[141], stage123[142], stage123[143], stage123[144], stage123[145]},
      {stage125[207], stage124[180], stage123[258], stage122[195], stage121[198]}
   );
   gpc615_5 gpc615_5_6060(
      {stage121[146], stage121[147], stage121[148], stage121[149], stage121[150]},
      {stage122[133]},
      {stage123[146], stage123[147], stage123[148], stage123[149], stage123[150], stage123[151]},
      {stage125[208], stage124[181], stage123[259], stage122[196], stage121[199]}
   );
   gpc615_5 gpc615_5_6061(
      {stage121[151], stage121[152], stage121[153], stage121[154], stage121[155]},
      {stage122[134]},
      {stage123[152], stage123[153], stage123[154], stage123[155], stage123[156], stage123[157]},
      {stage125[209], stage124[182], stage123[260], stage122[197], stage121[200]}
   );
   gpc615_5 gpc615_5_6062(
      {stage121[156], stage121[157], stage121[158], stage121[159], stage121[160]},
      {stage122[135]},
      {stage123[158], stage123[159], stage123[160], stage123[161], stage123[162], stage123[163]},
      {stage125[210], stage124[183], stage123[261], stage122[198], stage121[201]}
   );
   gpc615_5 gpc615_5_6063(
      {stage121[161], stage121[162], stage121[163], stage121[164], stage121[165]},
      {stage122[136]},
      {stage123[164], stage123[165], stage123[166], stage123[167], stage123[168], stage123[169]},
      {stage125[211], stage124[184], stage123[262], stage122[199], stage121[202]}
   );
   gpc615_5 gpc615_5_6064(
      {stage121[166], stage121[167], stage121[168], stage121[169], stage121[170]},
      {stage122[137]},
      {stage123[170], stage123[171], stage123[172], stage123[173], stage123[174], stage123[175]},
      {stage125[212], stage124[185], stage123[263], stage122[200], stage121[203]}
   );
   gpc615_5 gpc615_5_6065(
      {stage121[171], stage121[172], stage121[173], stage121[174], stage121[175]},
      {stage122[138]},
      {stage123[176], stage123[177], stage123[178], stage123[179], stage123[180], stage123[181]},
      {stage125[213], stage124[186], stage123[264], stage122[201], stage121[204]}
   );
   gpc1_1 gpc1_1_6066(
      {stage122[139]},
      {stage122[202]}
   );
   gpc1_1 gpc1_1_6067(
      {stage122[140]},
      {stage122[203]}
   );
   gpc1_1 gpc1_1_6068(
      {stage122[141]},
      {stage122[204]}
   );
   gpc1_1 gpc1_1_6069(
      {stage122[142]},
      {stage122[205]}
   );
   gpc1_1 gpc1_1_6070(
      {stage122[143]},
      {stage122[206]}
   );
   gpc1_1 gpc1_1_6071(
      {stage122[144]},
      {stage122[207]}
   );
   gpc1_1 gpc1_1_6072(
      {stage122[145]},
      {stage122[208]}
   );
   gpc1_1 gpc1_1_6073(
      {stage122[146]},
      {stage122[209]}
   );
   gpc1_1 gpc1_1_6074(
      {stage122[147]},
      {stage122[210]}
   );
   gpc1_1 gpc1_1_6075(
      {stage122[148]},
      {stage122[211]}
   );
   gpc1_1 gpc1_1_6076(
      {stage122[149]},
      {stage122[212]}
   );
   gpc1_1 gpc1_1_6077(
      {stage122[150]},
      {stage122[213]}
   );
   gpc1_1 gpc1_1_6078(
      {stage122[151]},
      {stage122[214]}
   );
   gpc615_5 gpc615_5_6079(
      {stage122[152], stage122[153], stage122[154], stage122[155], stage122[156]},
      {stage123[182]},
      {stage124[128], stage124[129], stage124[130], stage124[131], stage124[132], stage124[133]},
      {stage126[189], stage125[214], stage124[187], stage123[265], stage122[215]}
   );
   gpc615_5 gpc615_5_6080(
      {stage122[157], stage122[158], stage122[159], stage122[160], stage122[161]},
      {stage123[183]},
      {stage124[134], stage124[135], stage124[136], stage124[137], stage124[138], stage124[139]},
      {stage126[190], stage125[215], stage124[188], stage123[266], stage122[216]}
   );
   gpc615_5 gpc615_5_6081(
      {stage122[162], stage122[163], stage122[164], stage122[165], stage122[166]},
      {stage123[184]},
      {stage124[140], stage124[141], stage124[142], stage124[143], stage124[144], stage124[145]},
      {stage126[191], stage125[216], stage124[189], stage123[267], stage122[217]}
   );
   gpc615_5 gpc615_5_6082(
      {stage122[167], stage122[168], stage122[169], stage122[170], stage122[171]},
      {stage123[185]},
      {stage124[146], stage124[147], stage124[148], stage124[149], stage124[150], stage124[151]},
      {stage126[192], stage125[217], stage124[190], stage123[268], stage122[218]}
   );
   gpc615_5 gpc615_5_6083(
      {stage122[172], stage122[173], stage122[174], stage122[175], stage122[176]},
      {stage123[186]},
      {stage124[152], stage124[153], stage124[154], stage124[155], stage124[156], stage124[157]},
      {stage126[193], stage125[218], stage124[191], stage123[269], stage122[219]}
   );
   gpc615_5 gpc615_5_6084(
      {stage122[177], stage122[178], stage122[179], stage122[180], stage122[181]},
      {stage123[187]},
      {stage124[158], stage124[159], stage124[160], stage124[161], stage124[162], stage124[163]},
      {stage126[194], stage125[219], stage124[192], stage123[270], stage122[220]}
   );
   gpc615_5 gpc615_5_6085(
      {stage122[182], stage122[183], stage122[184], stage122[185], stage122[186]},
      {stage123[188]},
      {stage124[164], stage124[165], stage124[166], stage124[167], stage124[168], stage124[169]},
      {stage126[195], stage125[220], stage124[193], stage123[271], stage122[221]}
   );
   gpc606_5 gpc606_5_6086(
      {stage123[189], stage123[190], stage123[191], stage123[192], stage123[193], stage123[194]},
      {stage125[128], stage125[129], stage125[130], stage125[131], stage125[132], stage125[133]},
      {stage127[212], stage126[196], stage125[221], stage124[194], stage123[272]}
   );
   gpc606_5 gpc606_5_6087(
      {stage123[195], stage123[196], stage123[197], stage123[198], stage123[199], stage123[200]},
      {stage125[134], stage125[135], stage125[136], stage125[137], stage125[138], stage125[139]},
      {stage127[213], stage126[197], stage125[222], stage124[195], stage123[273]}
   );
   gpc606_5 gpc606_5_6088(
      {stage123[201], stage123[202], stage123[203], stage123[204], stage123[205], stage123[206]},
      {stage125[140], stage125[141], stage125[142], stage125[143], stage125[144], stage125[145]},
      {stage127[214], stage126[198], stage125[223], stage124[196], stage123[274]}
   );
   gpc207_4 gpc207_4_6089(
      {stage123[207], stage123[208], stage123[209], stage123[210], stage123[211], stage123[212], stage123[213]},
      {stage125[146], stage125[147]},
      {stage126[199], stage125[224], stage124[197], stage123[275]}
   );
   gpc207_4 gpc207_4_6090(
      {stage123[214], stage123[215], stage123[216], stage123[217], stage123[218], stage123[219], stage123[220]},
      {stage125[148], stage125[149]},
      {stage126[200], stage125[225], stage124[198], stage123[276]}
   );
   gpc207_4 gpc207_4_6091(
      {stage123[221], stage123[222], stage123[223], stage123[224], stage123[225], stage123[226], stage123[227]},
      {stage125[150], stage125[151]},
      {stage126[201], stage125[226], stage124[199], stage123[277]}
   );
   gpc207_4 gpc207_4_6092(
      {stage123[228], stage123[229], stage123[230], stage123[231], stage123[232], stage123[233], stage123[234]},
      {stage125[152], stage125[153]},
      {stage126[202], stage125[227], stage124[200], stage123[278]}
   );
   gpc207_4 gpc207_4_6093(
      {stage123[235], stage123[236], stage123[237], stage123[238], stage123[239], stage123[240], stage123[241]},
      {stage125[154], stage125[155]},
      {stage126[203], stage125[228], stage124[201], stage123[279]}
   );
   gpc207_4 gpc207_4_6094(
      {stage123[242], stage123[243], stage123[244], stage123[245], stage123[246], stage123[247], stage123[248]},
      {stage125[156], stage125[157]},
      {stage126[204], stage125[229], stage124[202], stage123[280]}
   );
   gpc207_4 gpc207_4_6095(
      {stage123[249], stage123[250], stage123[251], stage123[252], stage123[253], stage123[254], stage123[255]},
      {stage125[158], stage125[159]},
      {stage126[205], stage125[230], stage124[203], stage123[281]}
   );
   gpc1_1 gpc1_1_6096(
      {stage124[170]},
      {stage124[204]}
   );
   gpc1_1 gpc1_1_6097(
      {stage124[171]},
      {stage124[205]}
   );
   gpc1_1 gpc1_1_6098(
      {stage124[172]},
      {stage124[206]}
   );
   gpc1_1 gpc1_1_6099(
      {stage124[173]},
      {stage124[207]}
   );
   gpc1_1 gpc1_1_6100(
      {stage124[174]},
      {stage124[208]}
   );
   gpc1_1 gpc1_1_6101(
      {stage124[175]},
      {stage124[209]}
   );
   gpc1_1 gpc1_1_6102(
      {stage124[176]},
      {stage124[210]}
   );
   gpc1_1 gpc1_1_6103(
      {stage124[177]},
      {stage124[211]}
   );
   gpc615_5 gpc615_5_6104(
      {stage125[160], stage125[161], stage125[162], stage125[163], stage125[164]},
      {stage126[128]},
      {stage127[128], stage127[129], stage127[130], stage127[131], stage127[132], stage127[133]},
      {stage129[12], stage128[31], stage127[215], stage126[206], stage125[231]}
   );
   gpc615_5 gpc615_5_6105(
      {stage125[165], stage125[166], stage125[167], stage125[168], stage125[169]},
      {stage126[129]},
      {stage127[134], stage127[135], stage127[136], stage127[137], stage127[138], stage127[139]},
      {stage129[13], stage128[32], stage127[216], stage126[207], stage125[232]}
   );
   gpc615_5 gpc615_5_6106(
      {stage125[170], stage125[171], stage125[172], stage125[173], stage125[174]},
      {stage126[130]},
      {stage127[140], stage127[141], stage127[142], stage127[143], stage127[144], stage127[145]},
      {stage129[14], stage128[33], stage127[217], stage126[208], stage125[233]}
   );
   gpc615_5 gpc615_5_6107(
      {stage125[175], stage125[176], stage125[177], stage125[178], stage125[179]},
      {stage126[131]},
      {stage127[146], stage127[147], stage127[148], stage127[149], stage127[150], stage127[151]},
      {stage129[15], stage128[34], stage127[218], stage126[209], stage125[234]}
   );
   gpc615_5 gpc615_5_6108(
      {stage125[180], stage125[181], stage125[182], stage125[183], stage125[184]},
      {stage126[132]},
      {stage127[152], stage127[153], stage127[154], stage127[155], stage127[156], stage127[157]},
      {stage129[16], stage128[35], stage127[219], stage126[210], stage125[235]}
   );
   gpc615_5 gpc615_5_6109(
      {stage125[185], stage125[186], stage125[187], stage125[188], stage125[189]},
      {stage126[133]},
      {stage127[158], stage127[159], stage127[160], stage127[161], stage127[162], stage127[163]},
      {stage129[17], stage128[36], stage127[220], stage126[211], stage125[236]}
   );
   gpc615_5 gpc615_5_6110(
      {stage125[190], stage125[191], stage125[192], stage125[193], stage125[194]},
      {stage126[134]},
      {stage127[164], stage127[165], stage127[166], stage127[167], stage127[168], stage127[169]},
      {stage129[18], stage128[37], stage127[221], stage126[212], stage125[237]}
   );
   gpc615_5 gpc615_5_6111(
      {stage125[195], stage125[196], stage125[197], stage125[198], stage125[199]},
      {stage126[135]},
      {stage127[170], stage127[171], stage127[172], stage127[173], stage127[174], stage127[175]},
      {stage129[19], stage128[38], stage127[222], stage126[213], stage125[238]}
   );
   gpc615_5 gpc615_5_6112(
      {stage125[200], stage125[201], stage125[202], stage125[203], stage125[204]},
      {stage126[136]},
      {stage127[176], stage127[177], stage127[178], stage127[179], stage127[180], stage127[181]},
      {stage129[20], stage128[39], stage127[223], stage126[214], stage125[239]}
   );
   gpc615_5 gpc615_5_6113(
      {1'h0, 1'h0, 1'h0, 1'h0, 1'h0},
      {stage126[137]},
      {stage127[182], stage127[183], stage127[184], stage127[185], stage127[186], stage127[187]},
      {stage129[21], stage128[40], stage127[224], stage126[215], stage125[240]}
   );
   gpc1_1 gpc1_1_6114(
      {stage126[138]},
      {stage126[216]}
   );
   gpc1_1 gpc1_1_6115(
      {stage126[139]},
      {stage126[217]}
   );
   gpc1_1 gpc1_1_6116(
      {stage126[140]},
      {stage126[218]}
   );
   gpc1_1 gpc1_1_6117(
      {stage126[141]},
      {stage126[219]}
   );
   gpc1_1 gpc1_1_6118(
      {stage126[142]},
      {stage126[220]}
   );
   gpc1_1 gpc1_1_6119(
      {stage126[143]},
      {stage126[221]}
   );
   gpc1_1 gpc1_1_6120(
      {stage126[144]},
      {stage126[222]}
   );
   gpc1_1 gpc1_1_6121(
      {stage126[145]},
      {stage126[223]}
   );
   gpc1_1 gpc1_1_6122(
      {stage126[146]},
      {stage126[224]}
   );
   gpc1_1 gpc1_1_6123(
      {stage126[147]},
      {stage126[225]}
   );
   gpc1_1 gpc1_1_6124(
      {stage126[148]},
      {stage126[226]}
   );
   gpc1_1 gpc1_1_6125(
      {stage126[149]},
      {stage126[227]}
   );
   gpc1_1 gpc1_1_6126(
      {stage126[150]},
      {stage126[228]}
   );
   gpc1_1 gpc1_1_6127(
      {stage126[151]},
      {stage126[229]}
   );
   gpc1_1 gpc1_1_6128(
      {stage126[152]},
      {stage126[230]}
   );
   gpc1_1 gpc1_1_6129(
      {stage126[153]},
      {stage126[231]}
   );
   gpc1_1 gpc1_1_6130(
      {stage126[154]},
      {stage126[232]}
   );
   gpc1_1 gpc1_1_6131(
      {stage126[155]},
      {stage126[233]}
   );
   gpc1_1 gpc1_1_6132(
      {stage126[156]},
      {stage126[234]}
   );
   gpc1_1 gpc1_1_6133(
      {stage126[157]},
      {stage126[235]}
   );
   gpc1_1 gpc1_1_6134(
      {stage126[158]},
      {stage126[236]}
   );
   gpc606_5 gpc606_5_6135(
      {stage126[159], stage126[160], stage126[161], stage126[162], stage126[163], stage126[164]},
      {stage128[0], stage128[1], stage128[2], stage128[3], stage128[4], stage128[5]},
      {stage130[0], stage129[22], stage128[41], stage127[225], stage126[237]}
   );
   gpc606_5 gpc606_5_6136(
      {stage126[165], stage126[166], stage126[167], stage126[168], stage126[169], stage126[170]},
      {stage128[6], stage128[7], stage128[8], stage128[9], stage128[10], stage128[11]},
      {stage130[1], stage129[23], stage128[42], stage127[226], stage126[238]}
   );
   gpc606_5 gpc606_5_6137(
      {stage126[171], stage126[172], stage126[173], stage126[174], stage126[175], stage126[176]},
      {stage128[12], stage128[13], stage128[14], stage128[15], stage128[16], stage128[17]},
      {stage130[2], stage129[24], stage128[43], stage127[227], stage126[239]}
   );
   gpc606_5 gpc606_5_6138(
      {stage126[177], stage126[178], stage126[179], stage126[180], stage126[181], stage126[182]},
      {stage128[18], stage128[19], stage128[20], stage128[21], stage128[22], stage128[23]},
      {stage130[3], stage129[25], stage128[44], stage127[228], stage126[240]}
   );
   gpc606_5 gpc606_5_6139(
      {stage126[183], stage126[184], stage126[185], stage126[186], stage126[187], stage126[188]},
      {stage128[24], stage128[25], stage128[26], stage128[27], stage128[28], stage128[29]},
      {stage130[4], stage129[26], stage128[45], stage127[229], stage126[241]}
   );
   gpc1_1 gpc1_1_6140(
      {stage127[188]},
      {stage127[230]}
   );
   gpc1_1 gpc1_1_6141(
      {stage127[189]},
      {stage127[231]}
   );
   gpc1_1 gpc1_1_6142(
      {stage127[190]},
      {stage127[232]}
   );
   gpc1_1 gpc1_1_6143(
      {stage127[191]},
      {stage127[233]}
   );
   gpc1_1 gpc1_1_6144(
      {stage127[192]},
      {stage127[234]}
   );
   gpc1_1 gpc1_1_6145(
      {stage127[193]},
      {stage127[235]}
   );
   gpc1_1 gpc1_1_6146(
      {stage127[194]},
      {stage127[236]}
   );
   gpc1_1 gpc1_1_6147(
      {stage127[195]},
      {stage127[237]}
   );
   gpc1_1 gpc1_1_6148(
      {stage127[196]},
      {stage127[238]}
   );
   gpc1_1 gpc1_1_6149(
      {stage127[197]},
      {stage127[239]}
   );
   gpc1_1 gpc1_1_6150(
      {stage127[198]},
      {stage127[240]}
   );
   gpc1_1 gpc1_1_6151(
      {stage127[199]},
      {stage127[241]}
   );
   gpc1_1 gpc1_1_6152(
      {stage127[200]},
      {stage127[242]}
   );
   gpc1_1 gpc1_1_6153(
      {stage127[201]},
      {stage127[243]}
   );
   gpc1_1 gpc1_1_6154(
      {stage127[202]},
      {stage127[244]}
   );
   gpc1_1 gpc1_1_6155(
      {stage127[203]},
      {stage127[245]}
   );
   gpc1_1 gpc1_1_6156(
      {stage127[204]},
      {stage127[246]}
   );
   gpc1_1 gpc1_1_6157(
      {stage127[205]},
      {stage127[247]}
   );
   gpc1_1 gpc1_1_6158(
      {stage127[206]},
      {stage127[248]}
   );
   gpc1_1 gpc1_1_6159(
      {stage127[207]},
      {stage127[249]}
   );
   gpc1_1 gpc1_1_6160(
      {stage127[208]},
      {stage127[250]}
   );
   gpc1_1 gpc1_1_6161(
      {stage127[209]},
      {stage127[251]}
   );
   gpc1_1 gpc1_1_6162(
      {stage127[210]},
      {stage127[252]}
   );
   gpc1_1 gpc1_1_6163(
      {stage127[211]},
      {stage127[253]}
   );
   gpc1_1 gpc1_1_6164(
      {stage128[30]},
      {stage128[46]}
   );
   gpc1_1 gpc1_1_6165(
      {stage129[0]},
      {stage129[27]}
   );
   gpc1_1 gpc1_1_6166(
      {stage129[1]},
      {stage129[28]}
   );
   gpc1_1 gpc1_1_6167(
      {stage129[2]},
      {stage129[29]}
   );
   gpc1_1 gpc1_1_6168(
      {stage129[3]},
      {stage129[30]}
   );
   gpc1_1 gpc1_1_6169(
      {stage129[4]},
      {stage129[31]}
   );
   gpc1_1 gpc1_1_6170(
      {stage129[5]},
      {stage129[32]}
   );
   gpc1_1 gpc1_1_6171(
      {stage129[6]},
      {stage129[33]}
   );
   gpc1_1 gpc1_1_6172(
      {stage129[7]},
      {stage129[34]}
   );
   gpc1_1 gpc1_1_6173(
      {stage129[8]},
      {stage129[35]}
   );
   gpc1_1 gpc1_1_6174(
      {stage129[9]},
      {stage129[36]}
   );
   gpc1_1 gpc1_1_6175(
      {stage129[10]},
      {stage129[37]}
   );
   gpc1_1 gpc1_1_6176(
      {stage129[11]},
      {stage129[38]}
   );
   gpc1_1 gpc1_1_6177(
      {stage000[170]},
      {stage000[180]}
   );
   gpc1_1 gpc1_1_6178(
      {stage000[171]},
      {stage000[181]}
   );
   gpc1_1 gpc1_1_6179(
      {stage000[172]},
      {stage000[182]}
   );
   gpc1_1 gpc1_1_6180(
      {stage000[173]},
      {stage000[183]}
   );
   gpc1_1 gpc1_1_6181(
      {stage000[174]},
      {stage000[184]}
   );
   gpc615_5 gpc615_5_6182(
      {stage000[175], stage000[176], stage000[177], stage000[178], stage000[179]},
      {stage001[183]},
      {stage002[189], stage002[190], stage002[191], stage002[192], stage002[193], stage002[194]},
      {stage004[232], stage003[197], stage002[219], stage001[210], stage000[185]}
   );
   gpc1_1 gpc1_1_6183(
      {stage001[184]},
      {stage001[211]}
   );
   gpc1_1 gpc1_1_6184(
      {stage001[185]},
      {stage001[212]}
   );
   gpc1_1 gpc1_1_6185(
      {stage001[186]},
      {stage001[213]}
   );
   gpc606_5 gpc606_5_6186(
      {stage001[187], stage001[188], stage001[189], stage001[190], stage001[191], stage001[192]},
      {stage003[176], stage003[177], stage003[178], stage003[179], stage003[180], stage003[181]},
      {stage005[245], stage004[233], stage003[198], stage002[220], stage001[214]}
   );
   gpc606_5 gpc606_5_6187(
      {stage001[193], stage001[194], stage001[195], stage001[196], stage001[197], stage001[198]},
      {stage003[182], stage003[183], stage003[184], stage003[185], stage003[186], stage003[187]},
      {stage005[246], stage004[234], stage003[199], stage002[221], stage001[215]}
   );
   gpc606_5 gpc606_5_6188(
      {stage001[199], stage001[200], stage001[201], stage001[202], stage001[203], stage001[204]},
      {stage003[188], stage003[189], stage003[190], stage003[191], stage003[192], stage003[193]},
      {stage005[247], stage004[235], stage003[200], stage002[222], stage001[216]}
   );
   gpc135_4 gpc135_4_6189(
      {stage001[205], stage001[206], stage001[207], stage001[208], stage001[209]},
      {stage002[195], stage002[196], stage002[197]},
      {stage003[194]},
      {stage004[236], stage003[201], stage002[223], stage001[217]}
   );
   gpc1_1 gpc1_1_6190(
      {stage002[198]},
      {stage002[224]}
   );
   gpc1_1 gpc1_1_6191(
      {stage002[199]},
      {stage002[225]}
   );
   gpc1_1 gpc1_1_6192(
      {stage002[200]},
      {stage002[226]}
   );
   gpc1_1 gpc1_1_6193(
      {stage002[201]},
      {stage002[227]}
   );
   gpc1_1 gpc1_1_6194(
      {stage002[202]},
      {stage002[228]}
   );
   gpc1_1 gpc1_1_6195(
      {stage002[203]},
      {stage002[229]}
   );
   gpc1_1 gpc1_1_6196(
      {stage002[204]},
      {stage002[230]}
   );
   gpc1_1 gpc1_1_6197(
      {stage002[205]},
      {stage002[231]}
   );
   gpc1_1 gpc1_1_6198(
      {stage002[206]},
      {stage002[232]}
   );
   gpc606_5 gpc606_5_6199(
      {stage002[207], stage002[208], stage002[209], stage002[210], stage002[211], stage002[212]},
      {stage004[186], stage004[187], stage004[188], stage004[189], stage004[190], stage004[191]},
      {stage006[226], stage005[248], stage004[237], stage003[202], stage002[233]}
   );
   gpc606_5 gpc606_5_6200(
      {stage002[213], stage002[214], stage002[215], stage002[216], stage002[217], stage002[218]},
      {stage004[192], stage004[193], stage004[194], stage004[195], stage004[196], stage004[197]},
      {stage006[227], stage005[249], stage004[238], stage003[203], stage002[234]}
   );
   gpc1_1 gpc1_1_6201(
      {stage003[195]},
      {stage003[204]}
   );
   gpc1_1 gpc1_1_6202(
      {stage003[196]},
      {stage003[205]}
   );
   gpc1_1 gpc1_1_6203(
      {stage004[198]},
      {stage004[239]}
   );
   gpc1_1 gpc1_1_6204(
      {stage004[199]},
      {stage004[240]}
   );
   gpc1_1 gpc1_1_6205(
      {stage004[200]},
      {stage004[241]}
   );
   gpc1_1 gpc1_1_6206(
      {stage004[201]},
      {stage004[242]}
   );
   gpc1_1 gpc1_1_6207(
      {stage004[202]},
      {stage004[243]}
   );
   gpc1_1 gpc1_1_6208(
      {stage004[203]},
      {stage004[244]}
   );
   gpc1_1 gpc1_1_6209(
      {stage004[204]},
      {stage004[245]}
   );
   gpc1_1 gpc1_1_6210(
      {stage004[205]},
      {stage004[246]}
   );
   gpc606_5 gpc606_5_6211(
      {stage004[206], stage004[207], stage004[208], stage004[209], stage004[210], stage004[211]},
      {stage006[188], stage006[189], stage006[190], stage006[191], stage006[192], stage006[193]},
      {stage008[205], stage007[228], stage006[228], stage005[250], stage004[247]}
   );
   gpc615_5 gpc615_5_6212(
      {stage004[212], stage004[213], stage004[214], stage004[215], stage004[216]},
      {stage005[213]},
      {stage006[194], stage006[195], stage006[196], stage006[197], stage006[198], stage006[199]},
      {stage008[206], stage007[229], stage006[229], stage005[251], stage004[248]}
   );
   gpc615_5 gpc615_5_6213(
      {stage004[217], stage004[218], stage004[219], stage004[220], stage004[221]},
      {stage005[214]},
      {stage006[200], stage006[201], stage006[202], stage006[203], stage006[204], stage006[205]},
      {stage008[207], stage007[230], stage006[230], stage005[252], stage004[249]}
   );
   gpc615_5 gpc615_5_6214(
      {stage004[222], stage004[223], stage004[224], stage004[225], stage004[226]},
      {stage005[215]},
      {stage006[206], stage006[207], stage006[208], stage006[209], stage006[210], stage006[211]},
      {stage008[208], stage007[231], stage006[231], stage005[253], stage004[250]}
   );
   gpc615_5 gpc615_5_6215(
      {stage004[227], stage004[228], stage004[229], stage004[230], stage004[231]},
      {stage005[216]},
      {stage006[212], stage006[213], stage006[214], stage006[215], stage006[216], stage006[217]},
      {stage008[209], stage007[232], stage006[232], stage005[254], stage004[251]}
   );
   gpc1_1 gpc1_1_6216(
      {stage005[217]},
      {stage005[255]}
   );
   gpc1_1 gpc1_1_6217(
      {stage005[218]},
      {stage005[256]}
   );
   gpc1_1 gpc1_1_6218(
      {stage005[219]},
      {stage005[257]}
   );
   gpc1_1 gpc1_1_6219(
      {stage005[220]},
      {stage005[258]}
   );
   gpc606_5 gpc606_5_6220(
      {stage005[221], stage005[222], stage005[223], stage005[224], stage005[225], stage005[226]},
      {stage007[193], stage007[194], stage007[195], stage007[196], stage007[197], stage007[198]},
      {stage009[213], stage008[210], stage007[233], stage006[233], stage005[259]}
   );
   gpc606_5 gpc606_5_6221(
      {stage005[227], stage005[228], stage005[229], stage005[230], stage005[231], stage005[232]},
      {stage007[199], stage007[200], stage007[201], stage007[202], stage007[203], stage007[204]},
      {stage009[214], stage008[211], stage007[234], stage006[234], stage005[260]}
   );
   gpc606_5 gpc606_5_6222(
      {stage005[233], stage005[234], stage005[235], stage005[236], stage005[237], stage005[238]},
      {stage007[205], stage007[206], stage007[207], stage007[208], stage007[209], stage007[210]},
      {stage009[215], stage008[212], stage007[235], stage006[235], stage005[261]}
   );
   gpc606_5 gpc606_5_6223(
      {stage005[239], stage005[240], stage005[241], stage005[242], stage005[243], stage005[244]},
      {stage007[211], stage007[212], stage007[213], stage007[214], stage007[215], stage007[216]},
      {stage009[216], stage008[213], stage007[236], stage006[236], stage005[262]}
   );
   gpc1_1 gpc1_1_6224(
      {stage006[218]},
      {stage006[237]}
   );
   gpc1_1 gpc1_1_6225(
      {stage006[219]},
      {stage006[238]}
   );
   gpc1_1 gpc1_1_6226(
      {stage006[220]},
      {stage006[239]}
   );
   gpc1_1 gpc1_1_6227(
      {stage006[221]},
      {stage006[240]}
   );
   gpc1_1 gpc1_1_6228(
      {stage006[222]},
      {stage006[241]}
   );
   gpc1_1 gpc1_1_6229(
      {stage006[223]},
      {stage006[242]}
   );
   gpc1_1 gpc1_1_6230(
      {stage006[224]},
      {stage006[243]}
   );
   gpc1_1 gpc1_1_6231(
      {stage006[225]},
      {stage006[244]}
   );
   gpc1_1 gpc1_1_6232(
      {stage007[217]},
      {stage007[237]}
   );
   gpc1_1 gpc1_1_6233(
      {stage007[218]},
      {stage007[238]}
   );
   gpc1_1 gpc1_1_6234(
      {stage007[219]},
      {stage007[239]}
   );
   gpc1_1 gpc1_1_6235(
      {stage007[220]},
      {stage007[240]}
   );
   gpc1_1 gpc1_1_6236(
      {stage007[221]},
      {stage007[241]}
   );
   gpc1_1 gpc1_1_6237(
      {stage007[222]},
      {stage007[242]}
   );
   gpc615_5 gpc615_5_6238(
      {stage007[223], stage007[224], stage007[225], stage007[226], stage007[227]},
      {stage008[176]},
      {stage009[188], stage009[189], stage009[190], stage009[191], stage009[192], stage009[193]},
      {stage011[220], stage010[257], stage009[217], stage008[214], stage007[243]}
   );
   gpc1_1 gpc1_1_6239(
      {stage008[177]},
      {stage008[215]}
   );
   gpc1_1 gpc1_1_6240(
      {stage008[178]},
      {stage008[216]}
   );
   gpc1_1 gpc1_1_6241(
      {stage008[179]},
      {stage008[217]}
   );
   gpc1_1 gpc1_1_6242(
      {stage008[180]},
      {stage008[218]}
   );
   gpc606_5 gpc606_5_6243(
      {stage008[181], stage008[182], stage008[183], stage008[184], stage008[185], stage008[186]},
      {stage010[188], stage010[189], stage010[190], stage010[191], stage010[192], stage010[193]},
      {stage012[277], stage011[221], stage010[258], stage009[218], stage008[219]}
   );
   gpc606_5 gpc606_5_6244(
      {stage008[187], stage008[188], stage008[189], stage008[190], stage008[191], stage008[192]},
      {stage010[194], stage010[195], stage010[196], stage010[197], stage010[198], stage010[199]},
      {stage012[278], stage011[222], stage010[259], stage009[219], stage008[220]}
   );
   gpc606_5 gpc606_5_6245(
      {stage008[193], stage008[194], stage008[195], stage008[196], stage008[197], stage008[198]},
      {stage010[200], stage010[201], stage010[202], stage010[203], stage010[204], stage010[205]},
      {stage012[279], stage011[223], stage010[260], stage009[220], stage008[221]}
   );
   gpc606_5 gpc606_5_6246(
      {stage008[199], stage008[200], stage008[201], stage008[202], stage008[203], stage008[204]},
      {stage010[206], stage010[207], stage010[208], stage010[209], stage010[210], stage010[211]},
      {stage012[280], stage011[224], stage010[261], stage009[221], stage008[222]}
   );
   gpc1_1 gpc1_1_6247(
      {stage009[194]},
      {stage009[222]}
   );
   gpc1_1 gpc1_1_6248(
      {stage009[195]},
      {stage009[223]}
   );
   gpc1_1 gpc1_1_6249(
      {stage009[196]},
      {stage009[224]}
   );
   gpc1_1 gpc1_1_6250(
      {stage009[197]},
      {stage009[225]}
   );
   gpc1_1 gpc1_1_6251(
      {stage009[198]},
      {stage009[226]}
   );
   gpc1_1 gpc1_1_6252(
      {stage009[199]},
      {stage009[227]}
   );
   gpc1_1 gpc1_1_6253(
      {stage009[200]},
      {stage009[228]}
   );
   gpc606_5 gpc606_5_6254(
      {stage009[201], stage009[202], stage009[203], stage009[204], stage009[205], stage009[206]},
      {stage011[202], stage011[203], stage011[204], stage011[205], stage011[206], stage011[207]},
      {stage013[208], stage012[281], stage011[225], stage010[262], stage009[229]}
   );
   gpc606_5 gpc606_5_6255(
      {stage009[207], stage009[208], stage009[209], stage009[210], stage009[211], stage009[212]},
      {stage011[208], stage011[209], stage011[210], stage011[211], stage011[212], stage011[213]},
      {stage013[209], stage012[282], stage011[226], stage010[263], stage009[230]}
   );
   gpc1_1 gpc1_1_6256(
      {stage010[212]},
      {stage010[264]}
   );
   gpc1_1 gpc1_1_6257(
      {stage010[213]},
      {stage010[265]}
   );
   gpc1_1 gpc1_1_6258(
      {stage010[214]},
      {stage010[266]}
   );
   gpc1_1 gpc1_1_6259(
      {stage010[215]},
      {stage010[267]}
   );
   gpc1_1 gpc1_1_6260(
      {stage010[216]},
      {stage010[268]}
   );
   gpc1_1 gpc1_1_6261(
      {stage010[217]},
      {stage010[269]}
   );
   gpc1_1 gpc1_1_6262(
      {stage010[218]},
      {stage010[270]}
   );
   gpc1_1 gpc1_1_6263(
      {stage010[219]},
      {stage010[271]}
   );
   gpc1_1 gpc1_1_6264(
      {stage010[220]},
      {stage010[272]}
   );
   gpc606_5 gpc606_5_6265(
      {stage010[221], stage010[222], stage010[223], stage010[224], stage010[225], stage010[226]},
      {stage012[220], stage012[221], stage012[222], stage012[223], stage012[224], stage012[225]},
      {stage014[258], stage013[210], stage012[283], stage011[227], stage010[273]}
   );
   gpc606_5 gpc606_5_6266(
      {stage010[227], stage010[228], stage010[229], stage010[230], stage010[231], stage010[232]},
      {stage012[226], stage012[227], stage012[228], stage012[229], stage012[230], stage012[231]},
      {stage014[259], stage013[211], stage012[284], stage011[228], stage010[274]}
   );
   gpc606_5 gpc606_5_6267(
      {stage010[233], stage010[234], stage010[235], stage010[236], stage010[237], stage010[238]},
      {stage012[232], stage012[233], stage012[234], stage012[235], stage012[236], stage012[237]},
      {stage014[260], stage013[212], stage012[285], stage011[229], stage010[275]}
   );
   gpc606_5 gpc606_5_6268(
      {stage010[239], stage010[240], stage010[241], stage010[242], stage010[243], stage010[244]},
      {stage012[238], stage012[239], stage012[240], stage012[241], stage012[242], stage012[243]},
      {stage014[261], stage013[213], stage012[286], stage011[230], stage010[276]}
   );
   gpc606_5 gpc606_5_6269(
      {stage010[245], stage010[246], stage010[247], stage010[248], stage010[249], stage010[250]},
      {stage012[244], stage012[245], stage012[246], stage012[247], stage012[248], stage012[249]},
      {stage014[262], stage013[214], stage012[287], stage011[231], stage010[277]}
   );
   gpc606_5 gpc606_5_6270(
      {stage010[251], stage010[252], stage010[253], stage010[254], stage010[255], stage010[256]},
      {stage012[250], stage012[251], stage012[252], stage012[253], stage012[254], stage012[255]},
      {stage014[263], stage013[215], stage012[288], stage011[232], stage010[278]}
   );
   gpc1_1 gpc1_1_6271(
      {stage011[214]},
      {stage011[233]}
   );
   gpc1_1 gpc1_1_6272(
      {stage011[215]},
      {stage011[234]}
   );
   gpc1_1 gpc1_1_6273(
      {stage011[216]},
      {stage011[235]}
   );
   gpc1_1 gpc1_1_6274(
      {stage011[217]},
      {stage011[236]}
   );
   gpc1_1 gpc1_1_6275(
      {stage011[218]},
      {stage011[237]}
   );
   gpc1_1 gpc1_1_6276(
      {stage011[219]},
      {stage011[238]}
   );
   gpc1_1 gpc1_1_6277(
      {stage012[256]},
      {stage012[289]}
   );
   gpc1_1 gpc1_1_6278(
      {stage012[257]},
      {stage012[290]}
   );
   gpc1_1 gpc1_1_6279(
      {stage012[258]},
      {stage012[291]}
   );
   gpc1_1 gpc1_1_6280(
      {stage012[259]},
      {stage012[292]}
   );
   gpc1_1 gpc1_1_6281(
      {stage012[260]},
      {stage012[293]}
   );
   gpc1_1 gpc1_1_6282(
      {stage012[261]},
      {stage012[294]}
   );
   gpc1_1 gpc1_1_6283(
      {stage012[262]},
      {stage012[295]}
   );
   gpc1_1 gpc1_1_6284(
      {stage012[263]},
      {stage012[296]}
   );
   gpc1_1 gpc1_1_6285(
      {stage012[264]},
      {stage012[297]}
   );
   gpc1_1 gpc1_1_6286(
      {stage012[265]},
      {stage012[298]}
   );
   gpc1_1 gpc1_1_6287(
      {stage012[266]},
      {stage012[299]}
   );
   gpc1_1 gpc1_1_6288(
      {stage012[267]},
      {stage012[300]}
   );
   gpc1_1 gpc1_1_6289(
      {stage012[268]},
      {stage012[301]}
   );
   gpc1_1 gpc1_1_6290(
      {stage012[269]},
      {stage012[302]}
   );
   gpc1_1 gpc1_1_6291(
      {stage012[270]},
      {stage012[303]}
   );
   gpc1_1 gpc1_1_6292(
      {stage012[271]},
      {stage012[304]}
   );
   gpc1_1 gpc1_1_6293(
      {stage012[272]},
      {stage012[305]}
   );
   gpc1_1 gpc1_1_6294(
      {stage012[273]},
      {stage012[306]}
   );
   gpc1_1 gpc1_1_6295(
      {stage012[274]},
      {stage012[307]}
   );
   gpc1_1 gpc1_1_6296(
      {stage012[275]},
      {stage012[308]}
   );
   gpc1_1 gpc1_1_6297(
      {stage012[276]},
      {stage012[309]}
   );
   gpc1_1 gpc1_1_6298(
      {stage013[184]},
      {stage013[216]}
   );
   gpc1_1 gpc1_1_6299(
      {stage013[185]},
      {stage013[217]}
   );
   gpc1_1 gpc1_1_6300(
      {stage013[186]},
      {stage013[218]}
   );
   gpc1_1 gpc1_1_6301(
      {stage013[187]},
      {stage013[219]}
   );
   gpc1_1 gpc1_1_6302(
      {stage013[188]},
      {stage013[220]}
   );
   gpc1_1 gpc1_1_6303(
      {stage013[189]},
      {stage013[221]}
   );
   gpc1_1 gpc1_1_6304(
      {stage013[190]},
      {stage013[222]}
   );
   gpc1_1 gpc1_1_6305(
      {stage013[191]},
      {stage013[223]}
   );
   gpc1_1 gpc1_1_6306(
      {stage013[192]},
      {stage013[224]}
   );
   gpc1_1 gpc1_1_6307(
      {stage013[193]},
      {stage013[225]}
   );
   gpc1_1 gpc1_1_6308(
      {stage013[194]},
      {stage013[226]}
   );
   gpc1_1 gpc1_1_6309(
      {stage013[195]},
      {stage013[227]}
   );
   gpc1_1 gpc1_1_6310(
      {stage013[196]},
      {stage013[228]}
   );
   gpc1_1 gpc1_1_6311(
      {stage013[197]},
      {stage013[229]}
   );
   gpc1_1 gpc1_1_6312(
      {stage013[198]},
      {stage013[230]}
   );
   gpc1_1 gpc1_1_6313(
      {stage013[199]},
      {stage013[231]}
   );
   gpc1_1 gpc1_1_6314(
      {stage013[200]},
      {stage013[232]}
   );
   gpc1_1 gpc1_1_6315(
      {stage013[201]},
      {stage013[233]}
   );
   gpc606_5 gpc606_5_6316(
      {stage013[202], stage013[203], stage013[204], stage013[205], stage013[206], stage013[207]},
      {stage015[188], stage015[189], stage015[190], stage015[191], stage015[192], stage015[193]},
      {stage017[251], stage016[246], stage015[223], stage014[264], stage013[234]}
   );
   gpc1_1 gpc1_1_6317(
      {stage014[227]},
      {stage014[265]}
   );
   gpc1_1 gpc1_1_6318(
      {stage014[228]},
      {stage014[266]}
   );
   gpc1_1 gpc1_1_6319(
      {stage014[229]},
      {stage014[267]}
   );
   gpc1_1 gpc1_1_6320(
      {stage014[230]},
      {stage014[268]}
   );
   gpc1_1 gpc1_1_6321(
      {stage014[231]},
      {stage014[269]}
   );
   gpc1_1 gpc1_1_6322(
      {stage014[232]},
      {stage014[270]}
   );
   gpc1_1 gpc1_1_6323(
      {stage014[233]},
      {stage014[271]}
   );
   gpc1_1 gpc1_1_6324(
      {stage014[234]},
      {stage014[272]}
   );
   gpc1_1 gpc1_1_6325(
      {stage014[235]},
      {stage014[273]}
   );
   gpc1_1 gpc1_1_6326(
      {stage014[236]},
      {stage014[274]}
   );
   gpc1_1 gpc1_1_6327(
      {stage014[237]},
      {stage014[275]}
   );
   gpc1_1 gpc1_1_6328(
      {stage014[238]},
      {stage014[276]}
   );
   gpc1_1 gpc1_1_6329(
      {stage014[239]},
      {stage014[277]}
   );
   gpc1_1 gpc1_1_6330(
      {stage014[240]},
      {stage014[278]}
   );
   gpc1_1 gpc1_1_6331(
      {stage014[241]},
      {stage014[279]}
   );
   gpc1_1 gpc1_1_6332(
      {stage014[242]},
      {stage014[280]}
   );
   gpc1_1 gpc1_1_6333(
      {stage014[243]},
      {stage014[281]}
   );
   gpc1_1 gpc1_1_6334(
      {stage014[244]},
      {stage014[282]}
   );
   gpc1_1 gpc1_1_6335(
      {stage014[245]},
      {stage014[283]}
   );
   gpc1_1 gpc1_1_6336(
      {stage014[246]},
      {stage014[284]}
   );
   gpc1_1 gpc1_1_6337(
      {stage014[247]},
      {stage014[285]}
   );
   gpc615_5 gpc615_5_6338(
      {stage014[248], stage014[249], stage014[250], stage014[251], stage014[252]},
      {stage015[194]},
      {stage016[209], stage016[210], stage016[211], stage016[212], stage016[213], stage016[214]},
      {stage018[222], stage017[252], stage016[247], stage015[224], stage014[286]}
   );
   gpc615_5 gpc615_5_6339(
      {stage014[253], stage014[254], stage014[255], stage014[256], stage014[257]},
      {stage015[195]},
      {stage016[215], stage016[216], stage016[217], stage016[218], stage016[219], stage016[220]},
      {stage018[223], stage017[253], stage016[248], stage015[225], stage014[287]}
   );
   gpc1_1 gpc1_1_6340(
      {stage015[196]},
      {stage015[226]}
   );
   gpc1_1 gpc1_1_6341(
      {stage015[197]},
      {stage015[227]}
   );
   gpc1_1 gpc1_1_6342(
      {stage015[198]},
      {stage015[228]}
   );
   gpc1_1 gpc1_1_6343(
      {stage015[199]},
      {stage015[229]}
   );
   gpc1_1 gpc1_1_6344(
      {stage015[200]},
      {stage015[230]}
   );
   gpc1_1 gpc1_1_6345(
      {stage015[201]},
      {stage015[231]}
   );
   gpc1_1 gpc1_1_6346(
      {stage015[202]},
      {stage015[232]}
   );
   gpc1_1 gpc1_1_6347(
      {stage015[203]},
      {stage015[233]}
   );
   gpc1_1 gpc1_1_6348(
      {stage015[204]},
      {stage015[234]}
   );
   gpc1_1 gpc1_1_6349(
      {stage015[205]},
      {stage015[235]}
   );
   gpc1_1 gpc1_1_6350(
      {stage015[206]},
      {stage015[236]}
   );
   gpc606_5 gpc606_5_6351(
      {stage015[207], stage015[208], stage015[209], stage015[210], stage015[211], stage015[212]},
      {stage017[219], stage017[220], stage017[221], stage017[222], stage017[223], stage017[224]},
      {stage019[222], stage018[224], stage017[254], stage016[249], stage015[237]}
   );
   gpc615_5 gpc615_5_6352(
      {stage015[213], stage015[214], stage015[215], stage015[216], stage015[217]},
      {stage016[221]},
      {stage017[225], stage017[226], stage017[227], stage017[228], stage017[229], stage017[230]},
      {stage019[223], stage018[225], stage017[255], stage016[250], stage015[238]}
   );
   gpc615_5 gpc615_5_6353(
      {stage015[218], stage015[219], stage015[220], stage015[221], stage015[222]},
      {stage016[222]},
      {stage017[231], stage017[232], stage017[233], stage017[234], stage017[235], stage017[236]},
      {stage019[224], stage018[226], stage017[256], stage016[251], stage015[239]}
   );
   gpc1_1 gpc1_1_6354(
      {stage016[223]},
      {stage016[252]}
   );
   gpc1_1 gpc1_1_6355(
      {stage016[224]},
      {stage016[253]}
   );
   gpc1_1 gpc1_1_6356(
      {stage016[225]},
      {stage016[254]}
   );
   gpc1_1 gpc1_1_6357(
      {stage016[226]},
      {stage016[255]}
   );
   gpc1_1 gpc1_1_6358(
      {stage016[227]},
      {stage016[256]}
   );
   gpc1_1 gpc1_1_6359(
      {stage016[228]},
      {stage016[257]}
   );
   gpc1_1 gpc1_1_6360(
      {stage016[229]},
      {stage016[258]}
   );
   gpc1_1 gpc1_1_6361(
      {stage016[230]},
      {stage016[259]}
   );
   gpc1_1 gpc1_1_6362(
      {stage016[231]},
      {stage016[260]}
   );
   gpc1_1 gpc1_1_6363(
      {stage016[232]},
      {stage016[261]}
   );
   gpc1_1 gpc1_1_6364(
      {stage016[233]},
      {stage016[262]}
   );
   gpc1_1 gpc1_1_6365(
      {stage016[234]},
      {stage016[263]}
   );
   gpc1_1 gpc1_1_6366(
      {stage016[235]},
      {stage016[264]}
   );
   gpc1_1 gpc1_1_6367(
      {stage016[236]},
      {stage016[265]}
   );
   gpc1_1 gpc1_1_6368(
      {stage016[237]},
      {stage016[266]}
   );
   gpc1_1 gpc1_1_6369(
      {stage016[238]},
      {stage016[267]}
   );
   gpc1_1 gpc1_1_6370(
      {stage016[239]},
      {stage016[268]}
   );
   gpc1_1 gpc1_1_6371(
      {stage016[240]},
      {stage016[269]}
   );
   gpc1_1 gpc1_1_6372(
      {stage016[241]},
      {stage016[270]}
   );
   gpc1_1 gpc1_1_6373(
      {stage016[242]},
      {stage016[271]}
   );
   gpc1_1 gpc1_1_6374(
      {stage016[243]},
      {stage016[272]}
   );
   gpc1_1 gpc1_1_6375(
      {stage016[244]},
      {stage016[273]}
   );
   gpc1_1 gpc1_1_6376(
      {stage016[245]},
      {stage016[274]}
   );
   gpc1_1 gpc1_1_6377(
      {stage017[237]},
      {stage017[257]}
   );
   gpc1_1 gpc1_1_6378(
      {stage017[238]},
      {stage017[258]}
   );
   gpc1_1 gpc1_1_6379(
      {stage017[239]},
      {stage017[259]}
   );
   gpc1_1 gpc1_1_6380(
      {stage017[240]},
      {stage017[260]}
   );
   gpc1_1 gpc1_1_6381(
      {stage017[241]},
      {stage017[261]}
   );
   gpc1_1 gpc1_1_6382(
      {stage017[242]},
      {stage017[262]}
   );
   gpc1_1 gpc1_1_6383(
      {stage017[243]},
      {stage017[263]}
   );
   gpc1_1 gpc1_1_6384(
      {stage017[244]},
      {stage017[264]}
   );
   gpc606_5 gpc606_5_6385(
      {stage017[245], stage017[246], stage017[247], stage017[248], stage017[249], stage017[250]},
      {stage019[188], stage019[189], stage019[190], stage019[191], stage019[192], stage019[193]},
      {stage021[239], stage020[211], stage019[225], stage018[227], stage017[265]}
   );
   gpc1_1 gpc1_1_6386(
      {stage018[189]},
      {stage018[228]}
   );
   gpc1_1 gpc1_1_6387(
      {stage018[190]},
      {stage018[229]}
   );
   gpc1_1 gpc1_1_6388(
      {stage018[191]},
      {stage018[230]}
   );
   gpc1_1 gpc1_1_6389(
      {stage018[192]},
      {stage018[231]}
   );
   gpc1_1 gpc1_1_6390(
      {stage018[193]},
      {stage018[232]}
   );
   gpc1_1 gpc1_1_6391(
      {stage018[194]},
      {stage018[233]}
   );
   gpc1_1 gpc1_1_6392(
      {stage018[195]},
      {stage018[234]}
   );
   gpc1_1 gpc1_1_6393(
      {stage018[196]},
      {stage018[235]}
   );
   gpc1_1 gpc1_1_6394(
      {stage018[197]},
      {stage018[236]}
   );
   gpc606_5 gpc606_5_6395(
      {stage018[198], stage018[199], stage018[200], stage018[201], stage018[202], stage018[203]},
      {stage020[184], stage020[185], stage020[186], stage020[187], stage020[188], stage020[189]},
      {stage022[201], stage021[240], stage020[212], stage019[226], stage018[237]}
   );
   gpc606_5 gpc606_5_6396(
      {stage018[204], stage018[205], stage018[206], stage018[207], stage018[208], stage018[209]},
      {stage020[190], stage020[191], stage020[192], stage020[193], stage020[194], stage020[195]},
      {stage022[202], stage021[241], stage020[213], stage019[227], stage018[238]}
   );
   gpc606_5 gpc606_5_6397(
      {stage018[210], stage018[211], stage018[212], stage018[213], stage018[214], stage018[215]},
      {stage020[196], stage020[197], stage020[198], stage020[199], stage020[200], stage020[201]},
      {stage022[203], stage021[242], stage020[214], stage019[228], stage018[239]}
   );
   gpc606_5 gpc606_5_6398(
      {stage018[216], stage018[217], stage018[218], stage018[219], stage018[220], stage018[221]},
      {stage020[202], stage020[203], stage020[204], stage020[205], stage020[206], stage020[207]},
      {stage022[204], stage021[243], stage020[215], stage019[229], stage018[240]}
   );
   gpc1_1 gpc1_1_6399(
      {stage019[194]},
      {stage019[230]}
   );
   gpc1_1 gpc1_1_6400(
      {stage019[195]},
      {stage019[231]}
   );
   gpc1_1 gpc1_1_6401(
      {stage019[196]},
      {stage019[232]}
   );
   gpc1_1 gpc1_1_6402(
      {stage019[197]},
      {stage019[233]}
   );
   gpc1_1 gpc1_1_6403(
      {stage019[198]},
      {stage019[234]}
   );
   gpc1_1 gpc1_1_6404(
      {stage019[199]},
      {stage019[235]}
   );
   gpc1_1 gpc1_1_6405(
      {stage019[200]},
      {stage019[236]}
   );
   gpc1_1 gpc1_1_6406(
      {stage019[201]},
      {stage019[237]}
   );
   gpc1_1 gpc1_1_6407(
      {stage019[202]},
      {stage019[238]}
   );
   gpc1_1 gpc1_1_6408(
      {stage019[203]},
      {stage019[239]}
   );
   gpc1_1 gpc1_1_6409(
      {stage019[204]},
      {stage019[240]}
   );
   gpc1_1 gpc1_1_6410(
      {stage019[205]},
      {stage019[241]}
   );
   gpc1_1 gpc1_1_6411(
      {stage019[206]},
      {stage019[242]}
   );
   gpc615_5 gpc615_5_6412(
      {stage019[207], stage019[208], stage019[209], stage019[210], stage019[211]},
      {stage020[208]},
      {stage021[201], stage021[202], stage021[203], stage021[204], stage021[205], stage021[206]},
      {stage023[265], stage022[205], stage021[244], stage020[216], stage019[243]}
   );
   gpc1415_5 gpc1415_5_6413(
      {stage019[212], stage019[213], stage019[214], stage019[215], stage019[216]},
      {stage020[209]},
      {stage021[207], stage021[208], stage021[209], stage021[210]},
      {stage022[180]},
      {stage023[266], stage022[206], stage021[245], stage020[217], stage019[244]}
   );
   gpc1415_5 gpc1415_5_6414(
      {stage019[217], stage019[218], stage019[219], stage019[220], stage019[221]},
      {stage020[210]},
      {stage021[211], stage021[212], stage021[213], stage021[214]},
      {stage022[181]},
      {stage023[267], stage022[207], stage021[246], stage020[218], stage019[245]}
   );
   gpc1_1 gpc1_1_6415(
      {stage021[215]},
      {stage021[247]}
   );
   gpc1_1 gpc1_1_6416(
      {stage021[216]},
      {stage021[248]}
   );
   gpc1_1 gpc1_1_6417(
      {stage021[217]},
      {stage021[249]}
   );
   gpc1_1 gpc1_1_6418(
      {stage021[218]},
      {stage021[250]}
   );
   gpc1_1 gpc1_1_6419(
      {stage021[219]},
      {stage021[251]}
   );
   gpc1_1 gpc1_1_6420(
      {stage021[220]},
      {stage021[252]}
   );
   gpc1_1 gpc1_1_6421(
      {stage021[221]},
      {stage021[253]}
   );
   gpc1_1 gpc1_1_6422(
      {stage021[222]},
      {stage021[254]}
   );
   gpc1_1 gpc1_1_6423(
      {stage021[223]},
      {stage021[255]}
   );
   gpc1_1 gpc1_1_6424(
      {stage021[224]},
      {stage021[256]}
   );
   gpc1_1 gpc1_1_6425(
      {stage021[225]},
      {stage021[257]}
   );
   gpc1_1 gpc1_1_6426(
      {stage021[226]},
      {stage021[258]}
   );
   gpc1_1 gpc1_1_6427(
      {stage021[227]},
      {stage021[259]}
   );
   gpc1_1 gpc1_1_6428(
      {stage021[228]},
      {stage021[260]}
   );
   gpc1_1 gpc1_1_6429(
      {stage021[229]},
      {stage021[261]}
   );
   gpc1_1 gpc1_1_6430(
      {stage021[230]},
      {stage021[262]}
   );
   gpc1_1 gpc1_1_6431(
      {stage021[231]},
      {stage021[263]}
   );
   gpc1_1 gpc1_1_6432(
      {stage021[232]},
      {stage021[264]}
   );
   gpc1_1 gpc1_1_6433(
      {stage021[233]},
      {stage021[265]}
   );
   gpc1_1 gpc1_1_6434(
      {stage021[234]},
      {stage021[266]}
   );
   gpc1_1 gpc1_1_6435(
      {stage021[235]},
      {stage021[267]}
   );
   gpc1_1 gpc1_1_6436(
      {stage021[236]},
      {stage021[268]}
   );
   gpc1_1 gpc1_1_6437(
      {stage021[237]},
      {stage021[269]}
   );
   gpc1_1 gpc1_1_6438(
      {stage021[238]},
      {stage021[270]}
   );
   gpc1_1 gpc1_1_6439(
      {stage022[182]},
      {stage022[208]}
   );
   gpc1_1 gpc1_1_6440(
      {stage022[183]},
      {stage022[209]}
   );
   gpc1_1 gpc1_1_6441(
      {stage022[184]},
      {stage022[210]}
   );
   gpc1_1 gpc1_1_6442(
      {stage022[185]},
      {stage022[211]}
   );
   gpc615_5 gpc615_5_6443(
      {stage022[186], stage022[187], stage022[188], stage022[189], stage022[190]},
      {stage023[223]},
      {stage024[188], stage024[189], stage024[190], stage024[191], stage024[192], stage024[193]},
      {stage026[222], stage025[257], stage024[225], stage023[268], stage022[212]}
   );
   gpc615_5 gpc615_5_6444(
      {stage022[191], stage022[192], stage022[193], stage022[194], stage022[195]},
      {stage023[224]},
      {stage024[194], stage024[195], stage024[196], stage024[197], stage024[198], stage024[199]},
      {stage026[223], stage025[258], stage024[226], stage023[269], stage022[213]}
   );
   gpc615_5 gpc615_5_6445(
      {stage022[196], stage022[197], stage022[198], stage022[199], stage022[200]},
      {stage023[225]},
      {stage024[200], stage024[201], stage024[202], stage024[203], stage024[204], stage024[205]},
      {stage026[224], stage025[259], stage024[227], stage023[270], stage022[214]}
   );
   gpc1_1 gpc1_1_6446(
      {stage023[226]},
      {stage023[271]}
   );
   gpc1_1 gpc1_1_6447(
      {stage023[227]},
      {stage023[272]}
   );
   gpc1_1 gpc1_1_6448(
      {stage023[228]},
      {stage023[273]}
   );
   gpc1_1 gpc1_1_6449(
      {stage023[229]},
      {stage023[274]}
   );
   gpc1_1 gpc1_1_6450(
      {stage023[230]},
      {stage023[275]}
   );
   gpc1_1 gpc1_1_6451(
      {stage023[231]},
      {stage023[276]}
   );
   gpc1_1 gpc1_1_6452(
      {stage023[232]},
      {stage023[277]}
   );
   gpc1_1 gpc1_1_6453(
      {stage023[233]},
      {stage023[278]}
   );
   gpc1_1 gpc1_1_6454(
      {stage023[234]},
      {stage023[279]}
   );
   gpc1_1 gpc1_1_6455(
      {stage023[235]},
      {stage023[280]}
   );
   gpc1_1 gpc1_1_6456(
      {stage023[236]},
      {stage023[281]}
   );
   gpc1_1 gpc1_1_6457(
      {stage023[237]},
      {stage023[282]}
   );
   gpc1_1 gpc1_1_6458(
      {stage023[238]},
      {stage023[283]}
   );
   gpc1_1 gpc1_1_6459(
      {stage023[239]},
      {stage023[284]}
   );
   gpc1_1 gpc1_1_6460(
      {stage023[240]},
      {stage023[285]}
   );
   gpc1_1 gpc1_1_6461(
      {stage023[241]},
      {stage023[286]}
   );
   gpc1_1 gpc1_1_6462(
      {stage023[242]},
      {stage023[287]}
   );
   gpc1_1 gpc1_1_6463(
      {stage023[243]},
      {stage023[288]}
   );
   gpc1_1 gpc1_1_6464(
      {stage023[244]},
      {stage023[289]}
   );
   gpc1_1 gpc1_1_6465(
      {stage023[245]},
      {stage023[290]}
   );
   gpc1_1 gpc1_1_6466(
      {stage023[246]},
      {stage023[291]}
   );
   gpc606_5 gpc606_5_6467(
      {stage023[247], stage023[248], stage023[249], stage023[250], stage023[251], stage023[252]},
      {stage025[224], stage025[225], stage025[226], stage025[227], stage025[228], stage025[229]},
      {stage027[211], stage026[225], stage025[260], stage024[228], stage023[292]}
   );
   gpc606_5 gpc606_5_6468(
      {stage023[253], stage023[254], stage023[255], stage023[256], stage023[257], stage023[258]},
      {stage025[230], stage025[231], stage025[232], stage025[233], stage025[234], stage025[235]},
      {stage027[212], stage026[226], stage025[261], stage024[229], stage023[293]}
   );
   gpc606_5 gpc606_5_6469(
      {stage023[259], stage023[260], stage023[261], stage023[262], stage023[263], stage023[264]},
      {stage025[236], stage025[237], stage025[238], stage025[239], stage025[240], stage025[241]},
      {stage027[213], stage026[227], stage025[262], stage024[230], stage023[294]}
   );
   gpc1_1 gpc1_1_6470(
      {stage024[206]},
      {stage024[231]}
   );
   gpc1_1 gpc1_1_6471(
      {stage024[207]},
      {stage024[232]}
   );
   gpc1_1 gpc1_1_6472(
      {stage024[208]},
      {stage024[233]}
   );
   gpc1_1 gpc1_1_6473(
      {stage024[209]},
      {stage024[234]}
   );
   gpc1_1 gpc1_1_6474(
      {stage024[210]},
      {stage024[235]}
   );
   gpc1_1 gpc1_1_6475(
      {stage024[211]},
      {stage024[236]}
   );
   gpc1_1 gpc1_1_6476(
      {stage024[212]},
      {stage024[237]}
   );
   gpc1_1 gpc1_1_6477(
      {stage024[213]},
      {stage024[238]}
   );
   gpc1_1 gpc1_1_6478(
      {stage024[214]},
      {stage024[239]}
   );
   gpc1_1 gpc1_1_6479(
      {stage024[215]},
      {stage024[240]}
   );
   gpc1_1 gpc1_1_6480(
      {stage024[216]},
      {stage024[241]}
   );
   gpc1_1 gpc1_1_6481(
      {stage024[217]},
      {stage024[242]}
   );
   gpc1_1 gpc1_1_6482(
      {stage024[218]},
      {stage024[243]}
   );
   gpc606_5 gpc606_5_6483(
      {stage024[219], stage024[220], stage024[221], stage024[222], stage024[223], stage024[224]},
      {stage026[191], stage026[192], stage026[193], stage026[194], stage026[195], stage026[196]},
      {stage028[224], stage027[214], stage026[228], stage025[263], stage024[244]}
   );
   gpc1_1 gpc1_1_6484(
      {stage025[242]},
      {stage025[264]}
   );
   gpc1_1 gpc1_1_6485(
      {stage025[243]},
      {stage025[265]}
   );
   gpc1_1 gpc1_1_6486(
      {stage025[244]},
      {stage025[266]}
   );
   gpc1_1 gpc1_1_6487(
      {stage025[245]},
      {stage025[267]}
   );
   gpc1_1 gpc1_1_6488(
      {stage025[246]},
      {stage025[268]}
   );
   gpc1_1 gpc1_1_6489(
      {stage025[247]},
      {stage025[269]}
   );
   gpc1_1 gpc1_1_6490(
      {stage025[248]},
      {stage025[270]}
   );
   gpc1_1 gpc1_1_6491(
      {stage025[249]},
      {stage025[271]}
   );
   gpc1_1 gpc1_1_6492(
      {stage025[250]},
      {stage025[272]}
   );
   gpc1_1 gpc1_1_6493(
      {stage025[251]},
      {stage025[273]}
   );
   gpc1_1 gpc1_1_6494(
      {stage025[252]},
      {stage025[274]}
   );
   gpc1_1 gpc1_1_6495(
      {stage025[253]},
      {stage025[275]}
   );
   gpc1_1 gpc1_1_6496(
      {stage025[254]},
      {stage025[276]}
   );
   gpc1_1 gpc1_1_6497(
      {stage025[255]},
      {stage025[277]}
   );
   gpc1_1 gpc1_1_6498(
      {stage025[256]},
      {stage025[278]}
   );
   gpc1_1 gpc1_1_6499(
      {stage026[197]},
      {stage026[229]}
   );
   gpc606_5 gpc606_5_6500(
      {stage026[198], stage026[199], stage026[200], stage026[201], stage026[202], stage026[203]},
      {stage028[182], stage028[183], stage028[184], stage028[185], stage028[186], stage028[187]},
      {stage030[210], stage029[251], stage028[225], stage027[215], stage026[230]}
   );
   gpc606_5 gpc606_5_6501(
      {stage026[204], stage026[205], stage026[206], stage026[207], stage026[208], stage026[209]},
      {stage028[188], stage028[189], stage028[190], stage028[191], stage028[192], stage028[193]},
      {stage030[211], stage029[252], stage028[226], stage027[216], stage026[231]}
   );
   gpc606_5 gpc606_5_6502(
      {stage026[210], stage026[211], stage026[212], stage026[213], stage026[214], stage026[215]},
      {stage028[194], stage028[195], stage028[196], stage028[197], stage028[198], stage028[199]},
      {stage030[212], stage029[253], stage028[227], stage027[217], stage026[232]}
   );
   gpc606_5 gpc606_5_6503(
      {stage026[216], stage026[217], stage026[218], stage026[219], stage026[220], stage026[221]},
      {stage028[200], stage028[201], stage028[202], stage028[203], stage028[204], stage028[205]},
      {stage030[213], stage029[254], stage028[228], stage027[218], stage026[233]}
   );
   gpc1_1 gpc1_1_6504(
      {stage027[176]},
      {stage027[219]}
   );
   gpc1_1 gpc1_1_6505(
      {stage027[177]},
      {stage027[220]}
   );
   gpc1_1 gpc1_1_6506(
      {stage027[178]},
      {stage027[221]}
   );
   gpc1_1 gpc1_1_6507(
      {stage027[179]},
      {stage027[222]}
   );
   gpc1_1 gpc1_1_6508(
      {stage027[180]},
      {stage027[223]}
   );
   gpc606_5 gpc606_5_6509(
      {stage027[181], stage027[182], stage027[183], stage027[184], stage027[185], stage027[186]},
      {stage029[204], stage029[205], stage029[206], stage029[207], stage029[208], stage029[209]},
      {stage031[210], stage030[214], stage029[255], stage028[229], stage027[224]}
   );
   gpc606_5 gpc606_5_6510(
      {stage027[187], stage027[188], stage027[189], stage027[190], stage027[191], stage027[192]},
      {stage029[210], stage029[211], stage029[212], stage029[213], stage029[214], stage029[215]},
      {stage031[211], stage030[215], stage029[256], stage028[230], stage027[225]}
   );
   gpc606_5 gpc606_5_6511(
      {stage027[193], stage027[194], stage027[195], stage027[196], stage027[197], stage027[198]},
      {stage029[216], stage029[217], stage029[218], stage029[219], stage029[220], stage029[221]},
      {stage031[212], stage030[216], stage029[257], stage028[231], stage027[226]}
   );
   gpc606_5 gpc606_5_6512(
      {stage027[199], stage027[200], stage027[201], stage027[202], stage027[203], stage027[204]},
      {stage029[222], stage029[223], stage029[224], stage029[225], stage029[226], stage029[227]},
      {stage031[213], stage030[217], stage029[258], stage028[232], stage027[227]}
   );
   gpc606_5 gpc606_5_6513(
      {stage027[205], stage027[206], stage027[207], stage027[208], stage027[209], stage027[210]},
      {stage029[228], stage029[229], stage029[230], stage029[231], stage029[232], stage029[233]},
      {stage031[214], stage030[218], stage029[259], stage028[233], stage027[228]}
   );
   gpc1_1 gpc1_1_6514(
      {stage028[206]},
      {stage028[234]}
   );
   gpc1_1 gpc1_1_6515(
      {stage028[207]},
      {stage028[235]}
   );
   gpc606_5 gpc606_5_6516(
      {stage028[208], stage028[209], stage028[210], stage028[211], stage028[212], stage028[213]},
      {stage030[184], stage030[185], stage030[186], stage030[187], stage030[188], stage030[189]},
      {stage032[263], stage031[215], stage030[219], stage029[260], stage028[236]}
   );
   gpc615_5 gpc615_5_6517(
      {stage028[214], stage028[215], stage028[216], stage028[217], stage028[218]},
      {stage029[234]},
      {stage030[190], stage030[191], stage030[192], stage030[193], stage030[194], stage030[195]},
      {stage032[264], stage031[216], stage030[220], stage029[261], stage028[237]}
   );
   gpc615_5 gpc615_5_6518(
      {stage028[219], stage028[220], stage028[221], stage028[222], stage028[223]},
      {stage029[235]},
      {stage030[196], stage030[197], stage030[198], stage030[199], stage030[200], stage030[201]},
      {stage032[265], stage031[217], stage030[221], stage029[262], stage028[238]}
   );
   gpc1_1 gpc1_1_6519(
      {stage029[236]},
      {stage029[263]}
   );
   gpc1_1 gpc1_1_6520(
      {stage029[237]},
      {stage029[264]}
   );
   gpc1_1 gpc1_1_6521(
      {stage029[238]},
      {stage029[265]}
   );
   gpc1_1 gpc1_1_6522(
      {stage029[239]},
      {stage029[266]}
   );
   gpc1_1 gpc1_1_6523(
      {stage029[240]},
      {stage029[267]}
   );
   gpc1_1 gpc1_1_6524(
      {stage029[241]},
      {stage029[268]}
   );
   gpc1_1 gpc1_1_6525(
      {stage029[242]},
      {stage029[269]}
   );
   gpc1_1 gpc1_1_6526(
      {stage029[243]},
      {stage029[270]}
   );
   gpc1_1 gpc1_1_6527(
      {stage029[244]},
      {stage029[271]}
   );
   gpc1_1 gpc1_1_6528(
      {stage029[245]},
      {stage029[272]}
   );
   gpc615_5 gpc615_5_6529(
      {stage029[246], stage029[247], stage029[248], stage029[249], stage029[250]},
      {stage030[202]},
      {stage031[171], stage031[172], stage031[173], stage031[174], stage031[175], stage031[176]},
      {stage033[266], stage032[266], stage031[218], stage030[222], stage029[273]}
   );
   gpc1_1 gpc1_1_6530(
      {stage030[203]},
      {stage030[223]}
   );
   gpc1_1 gpc1_1_6531(
      {stage030[204]},
      {stage030[224]}
   );
   gpc1_1 gpc1_1_6532(
      {stage030[205]},
      {stage030[225]}
   );
   gpc1_1 gpc1_1_6533(
      {stage030[206]},
      {stage030[226]}
   );
   gpc1_1 gpc1_1_6534(
      {stage030[207]},
      {stage030[227]}
   );
   gpc1_1 gpc1_1_6535(
      {stage030[208]},
      {stage030[228]}
   );
   gpc1_1 gpc1_1_6536(
      {stage030[209]},
      {stage030[229]}
   );
   gpc1_1 gpc1_1_6537(
      {stage031[177]},
      {stage031[219]}
   );
   gpc1_1 gpc1_1_6538(
      {stage031[178]},
      {stage031[220]}
   );
   gpc1_1 gpc1_1_6539(
      {stage031[179]},
      {stage031[221]}
   );
   gpc1_1 gpc1_1_6540(
      {stage031[180]},
      {stage031[222]}
   );
   gpc1_1 gpc1_1_6541(
      {stage031[181]},
      {stage031[223]}
   );
   gpc1_1 gpc1_1_6542(
      {stage031[182]},
      {stage031[224]}
   );
   gpc1_1 gpc1_1_6543(
      {stage031[183]},
      {stage031[225]}
   );
   gpc1_1 gpc1_1_6544(
      {stage031[184]},
      {stage031[226]}
   );
   gpc1_1 gpc1_1_6545(
      {stage031[185]},
      {stage031[227]}
   );
   gpc1_1 gpc1_1_6546(
      {stage031[186]},
      {stage031[228]}
   );
   gpc1_1 gpc1_1_6547(
      {stage031[187]},
      {stage031[229]}
   );
   gpc1_1 gpc1_1_6548(
      {stage031[188]},
      {stage031[230]}
   );
   gpc1_1 gpc1_1_6549(
      {stage031[189]},
      {stage031[231]}
   );
   gpc1_1 gpc1_1_6550(
      {stage031[190]},
      {stage031[232]}
   );
   gpc1_1 gpc1_1_6551(
      {stage031[191]},
      {stage031[233]}
   );
   gpc615_5 gpc615_5_6552(
      {stage031[192], stage031[193], stage031[194], stage031[195], stage031[196]},
      {stage032[223]},
      {stage033[216], stage033[217], stage033[218], stage033[219], stage033[220], stage033[221]},
      {stage035[237], stage034[262], stage033[267], stage032[267], stage031[234]}
   );
   gpc615_5 gpc615_5_6553(
      {stage031[197], stage031[198], stage031[199], stage031[200], stage031[201]},
      {stage032[224]},
      {stage033[222], stage033[223], stage033[224], stage033[225], stage033[226], stage033[227]},
      {stage035[238], stage034[263], stage033[268], stage032[268], stage031[235]}
   );
   gpc615_5 gpc615_5_6554(
      {stage031[202], stage031[203], stage031[204], stage031[205], stage031[206]},
      {stage032[225]},
      {stage033[228], stage033[229], stage033[230], stage033[231], stage033[232], stage033[233]},
      {stage035[239], stage034[264], stage033[269], stage032[269], stage031[236]}
   );
   gpc1343_5 gpc1343_5_6555(
      {stage031[207], stage031[208], stage031[209]},
      {stage032[226], stage032[227], stage032[228], stage032[229]},
      {stage033[234], stage033[235], stage033[236]},
      {stage034[211]},
      {stage035[240], stage034[265], stage033[270], stage032[270], stage031[237]}
   );
   gpc1_1 gpc1_1_6556(
      {stage032[230]},
      {stage032[271]}
   );
   gpc1_1 gpc1_1_6557(
      {stage032[231]},
      {stage032[272]}
   );
   gpc1_1 gpc1_1_6558(
      {stage032[232]},
      {stage032[273]}
   );
   gpc1_1 gpc1_1_6559(
      {stage032[233]},
      {stage032[274]}
   );
   gpc1_1 gpc1_1_6560(
      {stage032[234]},
      {stage032[275]}
   );
   gpc1_1 gpc1_1_6561(
      {stage032[235]},
      {stage032[276]}
   );
   gpc1_1 gpc1_1_6562(
      {stage032[236]},
      {stage032[277]}
   );
   gpc1_1 gpc1_1_6563(
      {stage032[237]},
      {stage032[278]}
   );
   gpc1_1 gpc1_1_6564(
      {stage032[238]},
      {stage032[279]}
   );
   gpc606_5 gpc606_5_6565(
      {stage032[239], stage032[240], stage032[241], stage032[242], stage032[243], stage032[244]},
      {stage034[212], stage034[213], stage034[214], stage034[215], stage034[216], stage034[217]},
      {stage036[203], stage035[241], stage034[266], stage033[271], stage032[280]}
   );
   gpc606_5 gpc606_5_6566(
      {stage032[245], stage032[246], stage032[247], stage032[248], stage032[249], stage032[250]},
      {stage034[218], stage034[219], stage034[220], stage034[221], stage034[222], stage034[223]},
      {stage036[204], stage035[242], stage034[267], stage033[272], stage032[281]}
   );
   gpc606_5 gpc606_5_6567(
      {stage032[251], stage032[252], stage032[253], stage032[254], stage032[255], stage032[256]},
      {stage034[224], stage034[225], stage034[226], stage034[227], stage034[228], stage034[229]},
      {stage036[205], stage035[243], stage034[268], stage033[273], stage032[282]}
   );
   gpc606_5 gpc606_5_6568(
      {stage032[257], stage032[258], stage032[259], stage032[260], stage032[261], stage032[262]},
      {stage034[230], stage034[231], stage034[232], stage034[233], stage034[234], stage034[235]},
      {stage036[206], stage035[244], stage034[269], stage033[274], stage032[283]}
   );
   gpc1_1 gpc1_1_6569(
      {stage033[237]},
      {stage033[275]}
   );
   gpc1_1 gpc1_1_6570(
      {stage033[238]},
      {stage033[276]}
   );
   gpc1_1 gpc1_1_6571(
      {stage033[239]},
      {stage033[277]}
   );
   gpc1_1 gpc1_1_6572(
      {stage033[240]},
      {stage033[278]}
   );
   gpc1_1 gpc1_1_6573(
      {stage033[241]},
      {stage033[279]}
   );
   gpc606_5 gpc606_5_6574(
      {stage033[242], stage033[243], stage033[244], stage033[245], stage033[246], stage033[247]},
      {stage035[209], stage035[210], stage035[211], stage035[212], stage035[213], stage035[214]},
      {stage037[229], stage036[207], stage035[245], stage034[270], stage033[280]}
   );
   gpc606_5 gpc606_5_6575(
      {stage033[248], stage033[249], stage033[250], stage033[251], stage033[252], stage033[253]},
      {stage035[215], stage035[216], stage035[217], stage035[218], stage035[219], stage035[220]},
      {stage037[230], stage036[208], stage035[246], stage034[271], stage033[281]}
   );
   gpc606_5 gpc606_5_6576(
      {stage033[254], stage033[255], stage033[256], stage033[257], stage033[258], stage033[259]},
      {stage035[221], stage035[222], stage035[223], stage035[224], stage035[225], stage035[226]},
      {stage037[231], stage036[209], stage035[247], stage034[272], stage033[282]}
   );
   gpc606_5 gpc606_5_6577(
      {stage033[260], stage033[261], stage033[262], stage033[263], stage033[264], stage033[265]},
      {stage035[227], stage035[228], stage035[229], stage035[230], stage035[231], stage035[232]},
      {stage037[232], stage036[210], stage035[248], stage034[273], stage033[283]}
   );
   gpc1_1 gpc1_1_6578(
      {stage034[236]},
      {stage034[274]}
   );
   gpc615_5 gpc615_5_6579(
      {stage034[237], stage034[238], stage034[239], stage034[240], stage034[241]},
      {stage035[233]},
      {stage036[173], stage036[174], stage036[175], stage036[176], stage036[177], stage036[178]},
      {stage038[223], stage037[233], stage036[211], stage035[249], stage034[275]}
   );
   gpc615_5 gpc615_5_6580(
      {stage034[242], stage034[243], stage034[244], stage034[245], stage034[246]},
      {stage035[234]},
      {stage036[179], stage036[180], stage036[181], stage036[182], stage036[183], stage036[184]},
      {stage038[224], stage037[234], stage036[212], stage035[250], stage034[276]}
   );
   gpc615_5 gpc615_5_6581(
      {stage034[247], stage034[248], stage034[249], stage034[250], stage034[251]},
      {stage035[235]},
      {stage036[185], stage036[186], stage036[187], stage036[188], stage036[189], stage036[190]},
      {stage038[225], stage037[235], stage036[213], stage035[251], stage034[277]}
   );
   gpc615_5 gpc615_5_6582(
      {stage034[252], stage034[253], stage034[254], stage034[255], stage034[256]},
      {stage035[236]},
      {stage036[191], stage036[192], stage036[193], stage036[194], stage036[195], stage036[196]},
      {stage038[226], stage037[236], stage036[214], stage035[252], stage034[278]}
   );
   gpc615_5 gpc615_5_6583(
      {stage034[257], stage034[258], stage034[259], stage034[260], stage034[261]},
      {1'h0},
      {stage036[197], stage036[198], stage036[199], stage036[200], stage036[201], stage036[202]},
      {stage038[227], stage037[237], stage036[215], stage035[253], stage034[279]}
   );
   gpc1_1 gpc1_1_6584(
      {stage037[200]},
      {stage037[238]}
   );
   gpc1_1 gpc1_1_6585(
      {stage037[201]},
      {stage037[239]}
   );
   gpc1_1 gpc1_1_6586(
      {stage037[202]},
      {stage037[240]}
   );
   gpc1_1 gpc1_1_6587(
      {stage037[203]},
      {stage037[241]}
   );
   gpc1_1 gpc1_1_6588(
      {stage037[204]},
      {stage037[242]}
   );
   gpc1_1 gpc1_1_6589(
      {stage037[205]},
      {stage037[243]}
   );
   gpc1_1 gpc1_1_6590(
      {stage037[206]},
      {stage037[244]}
   );
   gpc1_1 gpc1_1_6591(
      {stage037[207]},
      {stage037[245]}
   );
   gpc1_1 gpc1_1_6592(
      {stage037[208]},
      {stage037[246]}
   );
   gpc1_1 gpc1_1_6593(
      {stage037[209]},
      {stage037[247]}
   );
   gpc1_1 gpc1_1_6594(
      {stage037[210]},
      {stage037[248]}
   );
   gpc1_1 gpc1_1_6595(
      {stage037[211]},
      {stage037[249]}
   );
   gpc1_1 gpc1_1_6596(
      {stage037[212]},
      {stage037[250]}
   );
   gpc1_1 gpc1_1_6597(
      {stage037[213]},
      {stage037[251]}
   );
   gpc1_1 gpc1_1_6598(
      {stage037[214]},
      {stage037[252]}
   );
   gpc1_1 gpc1_1_6599(
      {stage037[215]},
      {stage037[253]}
   );
   gpc1_1 gpc1_1_6600(
      {stage037[216]},
      {stage037[254]}
   );
   gpc1_1 gpc1_1_6601(
      {stage037[217]},
      {stage037[255]}
   );
   gpc1_1 gpc1_1_6602(
      {stage037[218]},
      {stage037[256]}
   );
   gpc2135_5 gpc2135_5_6603(
      {stage037[219], stage037[220], stage037[221], stage037[222], stage037[223]},
      {stage038[193], stage038[194], stage038[195]},
      {stage039[189]},
      {stage040[218], stage040[219]},
      {stage041[237], stage040[268], stage039[224], stage038[228], stage037[257]}
   );
   gpc2135_5 gpc2135_5_6604(
      {stage037[224], stage037[225], stage037[226], stage037[227], stage037[228]},
      {stage038[196], stage038[197], stage038[198]},
      {stage039[190]},
      {stage040[220], stage040[221]},
      {stage041[238], stage040[269], stage039[225], stage038[229], stage037[258]}
   );
   gpc606_5 gpc606_5_6605(
      {stage038[199], stage038[200], stage038[201], stage038[202], stage038[203], stage038[204]},
      {stage040[222], stage040[223], stage040[224], stage040[225], stage040[226], stage040[227]},
      {stage042[247], stage041[239], stage040[270], stage039[226], stage038[230]}
   );
   gpc606_5 gpc606_5_6606(
      {stage038[205], stage038[206], stage038[207], stage038[208], stage038[209], stage038[210]},
      {stage040[228], stage040[229], stage040[230], stage040[231], stage040[232], stage040[233]},
      {stage042[248], stage041[240], stage040[271], stage039[227], stage038[231]}
   );
   gpc606_5 gpc606_5_6607(
      {stage038[211], stage038[212], stage038[213], stage038[214], stage038[215], stage038[216]},
      {stage040[234], stage040[235], stage040[236], stage040[237], stage040[238], stage040[239]},
      {stage042[249], stage041[241], stage040[272], stage039[228], stage038[232]}
   );
   gpc606_5 gpc606_5_6608(
      {stage038[217], stage038[218], stage038[219], stage038[220], stage038[221], stage038[222]},
      {stage040[240], stage040[241], stage040[242], stage040[243], stage040[244], stage040[245]},
      {stage042[250], stage041[242], stage040[273], stage039[229], stage038[233]}
   );
   gpc1_1 gpc1_1_6609(
      {stage039[191]},
      {stage039[230]}
   );
   gpc1_1 gpc1_1_6610(
      {stage039[192]},
      {stage039[231]}
   );
   gpc1_1 gpc1_1_6611(
      {stage039[193]},
      {stage039[232]}
   );
   gpc1_1 gpc1_1_6612(
      {stage039[194]},
      {stage039[233]}
   );
   gpc1_1 gpc1_1_6613(
      {stage039[195]},
      {stage039[234]}
   );
   gpc1_1 gpc1_1_6614(
      {stage039[196]},
      {stage039[235]}
   );
   gpc1_1 gpc1_1_6615(
      {stage039[197]},
      {stage039[236]}
   );
   gpc1_1 gpc1_1_6616(
      {stage039[198]},
      {stage039[237]}
   );
   gpc615_5 gpc615_5_6617(
      {stage039[199], stage039[200], stage039[201], stage039[202], stage039[203]},
      {stage040[246]},
      {stage041[202], stage041[203], stage041[204], stage041[205], stage041[206], stage041[207]},
      {stage043[196], stage042[251], stage041[243], stage040[274], stage039[238]}
   );
   gpc615_5 gpc615_5_6618(
      {stage039[204], stage039[205], stage039[206], stage039[207], stage039[208]},
      {stage040[247]},
      {stage041[208], stage041[209], stage041[210], stage041[211], stage041[212], stage041[213]},
      {stage043[197], stage042[252], stage041[244], stage040[275], stage039[239]}
   );
   gpc615_5 gpc615_5_6619(
      {stage039[209], stage039[210], stage039[211], stage039[212], stage039[213]},
      {stage040[248]},
      {stage041[214], stage041[215], stage041[216], stage041[217], stage041[218], stage041[219]},
      {stage043[198], stage042[253], stage041[245], stage040[276], stage039[240]}
   );
   gpc615_5 gpc615_5_6620(
      {stage039[214], stage039[215], stage039[216], stage039[217], stage039[218]},
      {stage040[249]},
      {stage041[220], stage041[221], stage041[222], stage041[223], stage041[224], stage041[225]},
      {stage043[199], stage042[254], stage041[246], stage040[277], stage039[241]}
   );
   gpc615_5 gpc615_5_6621(
      {stage039[219], stage039[220], stage039[221], stage039[222], stage039[223]},
      {stage040[250]},
      {stage041[226], stage041[227], stage041[228], stage041[229], stage041[230], stage041[231]},
      {stage043[200], stage042[255], stage041[247], stage040[278], stage039[242]}
   );
   gpc1_1 gpc1_1_6622(
      {stage040[251]},
      {stage040[279]}
   );
   gpc1_1 gpc1_1_6623(
      {stage040[252]},
      {stage040[280]}
   );
   gpc1_1 gpc1_1_6624(
      {stage040[253]},
      {stage040[281]}
   );
   gpc1_1 gpc1_1_6625(
      {stage040[254]},
      {stage040[282]}
   );
   gpc1_1 gpc1_1_6626(
      {stage040[255]},
      {stage040[283]}
   );
   gpc606_5 gpc606_5_6627(
      {stage040[256], stage040[257], stage040[258], stage040[259], stage040[260], stage040[261]},
      {stage042[209], stage042[210], stage042[211], stage042[212], stage042[213], stage042[214]},
      {stage044[208], stage043[201], stage042[256], stage041[248], stage040[284]}
   );
   gpc606_5 gpc606_5_6628(
      {stage040[262], stage040[263], stage040[264], stage040[265], stage040[266], stage040[267]},
      {stage042[215], stage042[216], stage042[217], stage042[218], stage042[219], stage042[220]},
      {stage044[209], stage043[202], stage042[257], stage041[249], stage040[285]}
   );
   gpc1_1 gpc1_1_6629(
      {stage041[232]},
      {stage041[250]}
   );
   gpc1_1 gpc1_1_6630(
      {stage041[233]},
      {stage041[251]}
   );
   gpc623_5 gpc623_5_6631(
      {stage041[234], stage041[235], stage041[236]},
      {stage042[221], stage042[222]},
      {stage043[166], stage043[167], stage043[168], stage043[169], stage043[170], stage043[171]},
      {stage045[250], stage044[210], stage043[203], stage042[258], stage041[252]}
   );
   gpc1_1 gpc1_1_6632(
      {stage042[223]},
      {stage042[259]}
   );
   gpc1_1 gpc1_1_6633(
      {stage042[224]},
      {stage042[260]}
   );
   gpc1_1 gpc1_1_6634(
      {stage042[225]},
      {stage042[261]}
   );
   gpc1_1 gpc1_1_6635(
      {stage042[226]},
      {stage042[262]}
   );
   gpc1_1 gpc1_1_6636(
      {stage042[227]},
      {stage042[263]}
   );
   gpc1_1 gpc1_1_6637(
      {stage042[228]},
      {stage042[264]}
   );
   gpc1_1 gpc1_1_6638(
      {stage042[229]},
      {stage042[265]}
   );
   gpc1_1 gpc1_1_6639(
      {stage042[230]},
      {stage042[266]}
   );
   gpc1_1 gpc1_1_6640(
      {stage042[231]},
      {stage042[267]}
   );
   gpc1_1 gpc1_1_6641(
      {stage042[232]},
      {stage042[268]}
   );
   gpc1_1 gpc1_1_6642(
      {stage042[233]},
      {stage042[269]}
   );
   gpc1_1 gpc1_1_6643(
      {stage042[234]},
      {stage042[270]}
   );
   gpc1_1 gpc1_1_6644(
      {stage042[235]},
      {stage042[271]}
   );
   gpc1_1 gpc1_1_6645(
      {stage042[236]},
      {stage042[272]}
   );
   gpc1_1 gpc1_1_6646(
      {stage042[237]},
      {stage042[273]}
   );
   gpc1_1 gpc1_1_6647(
      {stage042[238]},
      {stage042[274]}
   );
   gpc1_1 gpc1_1_6648(
      {stage042[239]},
      {stage042[275]}
   );
   gpc1_1 gpc1_1_6649(
      {stage042[240]},
      {stage042[276]}
   );
   gpc1_1 gpc1_1_6650(
      {stage042[241]},
      {stage042[277]}
   );
   gpc615_5 gpc615_5_6651(
      {stage042[242], stage042[243], stage042[244], stage042[245], stage042[246]},
      {stage043[172]},
      {stage044[179], stage044[180], stage044[181], stage044[182], stage044[183], stage044[184]},
      {stage046[249], stage045[251], stage044[211], stage043[204], stage042[278]}
   );
   gpc615_5 gpc615_5_6652(
      {stage043[173], stage043[174], stage043[175], stage043[176], stage043[177]},
      {stage044[185]},
      {stage045[204], stage045[205], stage045[206], stage045[207], stage045[208], stage045[209]},
      {stage047[198], stage046[250], stage045[252], stage044[212], stage043[205]}
   );
   gpc615_5 gpc615_5_6653(
      {stage043[178], stage043[179], stage043[180], stage043[181], stage043[182]},
      {stage044[186]},
      {stage045[210], stage045[211], stage045[212], stage045[213], stage045[214], stage045[215]},
      {stage047[199], stage046[251], stage045[253], stage044[213], stage043[206]}
   );
   gpc615_5 gpc615_5_6654(
      {stage043[183], stage043[184], stage043[185], stage043[186], stage043[187]},
      {stage044[187]},
      {stage045[216], stage045[217], stage045[218], stage045[219], stage045[220], stage045[221]},
      {stage047[200], stage046[252], stage045[254], stage044[214], stage043[207]}
   );
   gpc615_5 gpc615_5_6655(
      {stage043[188], stage043[189], stage043[190], stage043[191], stage043[192]},
      {stage044[188]},
      {stage045[222], stage045[223], stage045[224], stage045[225], stage045[226], stage045[227]},
      {stage047[201], stage046[253], stage045[255], stage044[215], stage043[208]}
   );
   gpc615_5 gpc615_5_6656(
      {stage043[193], stage043[194], stage043[195], 1'h0, 1'h0},
      {stage044[189]},
      {stage045[228], stage045[229], stage045[230], stage045[231], stage045[232], stage045[233]},
      {stage047[202], stage046[254], stage045[256], stage044[216], stage043[209]}
   );
   gpc606_5 gpc606_5_6657(
      {stage044[190], stage044[191], stage044[192], stage044[193], stage044[194], stage044[195]},
      {stage046[216], stage046[217], stage046[218], stage046[219], stage046[220], stage046[221]},
      {stage048[295], stage047[203], stage046[255], stage045[257], stage044[217]}
   );
   gpc606_5 gpc606_5_6658(
      {stage044[196], stage044[197], stage044[198], stage044[199], stage044[200], stage044[201]},
      {stage046[222], stage046[223], stage046[224], stage046[225], stage046[226], stage046[227]},
      {stage048[296], stage047[204], stage046[256], stage045[258], stage044[218]}
   );
   gpc606_5 gpc606_5_6659(
      {stage044[202], stage044[203], stage044[204], stage044[205], stage044[206], stage044[207]},
      {stage046[228], stage046[229], stage046[230], stage046[231], stage046[232], stage046[233]},
      {stage048[297], stage047[205], stage046[257], stage045[259], stage044[219]}
   );
   gpc1_1 gpc1_1_6660(
      {stage045[234]},
      {stage045[260]}
   );
   gpc1_1 gpc1_1_6661(
      {stage045[235]},
      {stage045[261]}
   );
   gpc1_1 gpc1_1_6662(
      {stage045[236]},
      {stage045[262]}
   );
   gpc1_1 gpc1_1_6663(
      {stage045[237]},
      {stage045[263]}
   );
   gpc606_5 gpc606_5_6664(
      {stage045[238], stage045[239], stage045[240], stage045[241], stage045[242], stage045[243]},
      {stage047[170], stage047[171], stage047[172], stage047[173], stage047[174], stage047[175]},
      {stage049[230], stage048[298], stage047[206], stage046[258], stage045[264]}
   );
   gpc606_5 gpc606_5_6665(
      {stage045[244], stage045[245], stage045[246], stage045[247], stage045[248], stage045[249]},
      {stage047[176], stage047[177], stage047[178], stage047[179], stage047[180], stage047[181]},
      {stage049[231], stage048[299], stage047[207], stage046[259], stage045[265]}
   );
   gpc615_5 gpc615_5_6666(
      {stage046[234], stage046[235], stage046[236], stage046[237], stage046[238]},
      {stage047[182]},
      {stage048[230], stage048[231], stage048[232], stage048[233], stage048[234], stage048[235]},
      {stage050[255], stage049[232], stage048[300], stage047[208], stage046[260]}
   );
   gpc615_5 gpc615_5_6667(
      {stage046[239], stage046[240], stage046[241], stage046[242], stage046[243]},
      {stage047[183]},
      {stage048[236], stage048[237], stage048[238], stage048[239], stage048[240], stage048[241]},
      {stage050[256], stage049[233], stage048[301], stage047[209], stage046[261]}
   );
   gpc615_5 gpc615_5_6668(
      {stage046[244], stage046[245], stage046[246], stage046[247], stage046[248]},
      {stage047[184]},
      {stage048[242], stage048[243], stage048[244], stage048[245], stage048[246], stage048[247]},
      {stage050[257], stage049[234], stage048[302], stage047[210], stage046[262]}
   );
   gpc1_1 gpc1_1_6669(
      {stage047[185]},
      {stage047[211]}
   );
   gpc1_1 gpc1_1_6670(
      {stage047[186]},
      {stage047[212]}
   );
   gpc1_1 gpc1_1_6671(
      {stage047[187]},
      {stage047[213]}
   );
   gpc1_1 gpc1_1_6672(
      {stage047[188]},
      {stage047[214]}
   );
   gpc1_1 gpc1_1_6673(
      {stage047[189]},
      {stage047[215]}
   );
   gpc1_1 gpc1_1_6674(
      {stage047[190]},
      {stage047[216]}
   );
   gpc1_1 gpc1_1_6675(
      {stage047[191]},
      {stage047[217]}
   );
   gpc1_1 gpc1_1_6676(
      {stage047[192]},
      {stage047[218]}
   );
   gpc1_1 gpc1_1_6677(
      {stage047[193]},
      {stage047[219]}
   );
   gpc1_1 gpc1_1_6678(
      {stage047[194]},
      {stage047[220]}
   );
   gpc1_1 gpc1_1_6679(
      {stage047[195]},
      {stage047[221]}
   );
   gpc1_1 gpc1_1_6680(
      {stage047[196]},
      {stage047[222]}
   );
   gpc1_1 gpc1_1_6681(
      {stage047[197]},
      {stage047[223]}
   );
   gpc1_1 gpc1_1_6682(
      {stage048[248]},
      {stage048[303]}
   );
   gpc1_1 gpc1_1_6683(
      {stage048[249]},
      {stage048[304]}
   );
   gpc1_1 gpc1_1_6684(
      {stage048[250]},
      {stage048[305]}
   );
   gpc1_1 gpc1_1_6685(
      {stage048[251]},
      {stage048[306]}
   );
   gpc1_1 gpc1_1_6686(
      {stage048[252]},
      {stage048[307]}
   );
   gpc1_1 gpc1_1_6687(
      {stage048[253]},
      {stage048[308]}
   );
   gpc1_1 gpc1_1_6688(
      {stage048[254]},
      {stage048[309]}
   );
   gpc1_1 gpc1_1_6689(
      {stage048[255]},
      {stage048[310]}
   );
   gpc1_1 gpc1_1_6690(
      {stage048[256]},
      {stage048[311]}
   );
   gpc1_1 gpc1_1_6691(
      {stage048[257]},
      {stage048[312]}
   );
   gpc1_1 gpc1_1_6692(
      {stage048[258]},
      {stage048[313]}
   );
   gpc1_1 gpc1_1_6693(
      {stage048[259]},
      {stage048[314]}
   );
   gpc606_5 gpc606_5_6694(
      {stage048[260], stage048[261], stage048[262], stage048[263], stage048[264], stage048[265]},
      {stage050[224], stage050[225], stage050[226], stage050[227], stage050[228], stage050[229]},
      {stage052[243], stage051[222], stage050[258], stage049[235], stage048[315]}
   );
   gpc606_5 gpc606_5_6695(
      {stage048[266], stage048[267], stage048[268], stage048[269], stage048[270], stage048[271]},
      {stage050[230], stage050[231], stage050[232], stage050[233], stage050[234], stage050[235]},
      {stage052[244], stage051[223], stage050[259], stage049[236], stage048[316]}
   );
   gpc606_5 gpc606_5_6696(
      {stage048[272], stage048[273], stage048[274], stage048[275], stage048[276], stage048[277]},
      {stage050[236], stage050[237], stage050[238], stage050[239], stage050[240], stage050[241]},
      {stage052[245], stage051[224], stage050[260], stage049[237], stage048[317]}
   );
   gpc606_5 gpc606_5_6697(
      {stage048[278], stage048[279], stage048[280], stage048[281], stage048[282], stage048[283]},
      {stage050[242], stage050[243], stage050[244], stage050[245], stage050[246], stage050[247]},
      {stage052[246], stage051[225], stage050[261], stage049[238], stage048[318]}
   );
   gpc606_5 gpc606_5_6698(
      {stage048[284], stage048[285], stage048[286], stage048[287], stage048[288], stage048[289]},
      {stage050[248], stage050[249], stage050[250], stage050[251], stage050[252], stage050[253]},
      {stage052[247], stage051[226], stage050[262], stage049[239], stage048[319]}
   );
   gpc1325_5 gpc1325_5_6699(
      {stage048[290], stage048[291], stage048[292], stage048[293], stage048[294]},
      {stage049[204], stage049[205]},
      {stage050[254], 1'h0, 1'h0},
      {stage051[167]},
      {stage052[248], stage051[227], stage050[263], stage049[240], stage048[320]}
   );
   gpc606_5 gpc606_5_6700(
      {stage049[206], stage049[207], stage049[208], stage049[209], stage049[210], stage049[211]},
      {stage051[168], stage051[169], stage051[170], stage051[171], stage051[172], stage051[173]},
      {stage053[212], stage052[249], stage051[228], stage050[264], stage049[241]}
   );
   gpc606_5 gpc606_5_6701(
      {stage049[212], stage049[213], stage049[214], stage049[215], stage049[216], stage049[217]},
      {stage051[174], stage051[175], stage051[176], stage051[177], stage051[178], stage051[179]},
      {stage053[213], stage052[250], stage051[229], stage050[265], stage049[242]}
   );
   gpc606_5 gpc606_5_6702(
      {stage049[218], stage049[219], stage049[220], stage049[221], stage049[222], stage049[223]},
      {stage051[180], stage051[181], stage051[182], stage051[183], stage051[184], stage051[185]},
      {stage053[214], stage052[251], stage051[230], stage050[266], stage049[243]}
   );
   gpc606_5 gpc606_5_6703(
      {stage049[224], stage049[225], stage049[226], stage049[227], stage049[228], stage049[229]},
      {stage051[186], stage051[187], stage051[188], stage051[189], stage051[190], stage051[191]},
      {stage053[215], stage052[252], stage051[231], stage050[267], stage049[244]}
   );
   gpc606_5 gpc606_5_6704(
      {stage051[192], stage051[193], stage051[194], stage051[195], stage051[196], stage051[197]},
      {stage053[171], stage053[172], stage053[173], stage053[174], stage053[175], stage053[176]},
      {stage055[247], stage054[234], stage053[216], stage052[253], stage051[232]}
   );
   gpc606_5 gpc606_5_6705(
      {stage051[198], stage051[199], stage051[200], stage051[201], stage051[202], stage051[203]},
      {stage053[177], stage053[178], stage053[179], stage053[180], stage053[181], stage053[182]},
      {stage055[248], stage054[235], stage053[217], stage052[254], stage051[233]}
   );
   gpc606_5 gpc606_5_6706(
      {stage051[204], stage051[205], stage051[206], stage051[207], stage051[208], stage051[209]},
      {stage053[183], stage053[184], stage053[185], stage053[186], stage053[187], stage053[188]},
      {stage055[249], stage054[236], stage053[218], stage052[255], stage051[234]}
   );
   gpc606_5 gpc606_5_6707(
      {stage051[210], stage051[211], stage051[212], stage051[213], stage051[214], stage051[215]},
      {stage053[189], stage053[190], stage053[191], stage053[192], stage053[193], stage053[194]},
      {stage055[250], stage054[237], stage053[219], stage052[256], stage051[235]}
   );
   gpc606_5 gpc606_5_6708(
      {stage051[216], stage051[217], stage051[218], stage051[219], stage051[220], stage051[221]},
      {stage053[195], stage053[196], stage053[197], stage053[198], stage053[199], stage053[200]},
      {stage055[251], stage054[238], stage053[220], stage052[257], stage051[236]}
   );
   gpc606_5 gpc606_5_6709(
      {stage052[214], stage052[215], stage052[216], stage052[217], stage052[218], stage052[219]},
      {stage054[205], stage054[206], stage054[207], stage054[208], stage054[209], stage054[210]},
      {stage056[235], stage055[252], stage054[239], stage053[221], stage052[258]}
   );
   gpc606_5 gpc606_5_6710(
      {stage052[220], stage052[221], stage052[222], stage052[223], stage052[224], stage052[225]},
      {stage054[211], stage054[212], stage054[213], stage054[214], stage054[215], stage054[216]},
      {stage056[236], stage055[253], stage054[240], stage053[222], stage052[259]}
   );
   gpc606_5 gpc606_5_6711(
      {stage052[226], stage052[227], stage052[228], stage052[229], stage052[230], stage052[231]},
      {stage054[217], stage054[218], stage054[219], stage054[220], stage054[221], stage054[222]},
      {stage056[237], stage055[254], stage054[241], stage053[223], stage052[260]}
   );
   gpc606_5 gpc606_5_6712(
      {stage052[232], stage052[233], stage052[234], stage052[235], stage052[236], stage052[237]},
      {stage054[223], stage054[224], stage054[225], stage054[226], stage054[227], stage054[228]},
      {stage056[238], stage055[255], stage054[242], stage053[224], stage052[261]}
   );
   gpc606_5 gpc606_5_6713(
      {stage052[238], stage052[239], stage052[240], stage052[241], stage052[242], 1'h0},
      {stage054[229], stage054[230], stage054[231], stage054[232], stage054[233], 1'h0},
      {stage056[239], stage055[256], stage054[243], stage053[225], stage052[262]}
   );
   gpc1_1 gpc1_1_6714(
      {stage053[201]},
      {stage053[226]}
   );
   gpc1_1 gpc1_1_6715(
      {stage053[202]},
      {stage053[227]}
   );
   gpc1_1 gpc1_1_6716(
      {stage053[203]},
      {stage053[228]}
   );
   gpc1_1 gpc1_1_6717(
      {stage053[204]},
      {stage053[229]}
   );
   gpc1_1 gpc1_1_6718(
      {stage053[205]},
      {stage053[230]}
   );
   gpc606_5 gpc606_5_6719(
      {stage053[206], stage053[207], stage053[208], stage053[209], stage053[210], stage053[211]},
      {stage055[199], stage055[200], stage055[201], stage055[202], stage055[203], stage055[204]},
      {stage057[233], stage056[240], stage055[257], stage054[244], stage053[231]}
   );
   gpc606_5 gpc606_5_6720(
      {stage055[205], stage055[206], stage055[207], stage055[208], stage055[209], stage055[210]},
      {stage057[184], stage057[185], stage057[186], stage057[187], stage057[188], stage057[189]},
      {stage059[267], stage058[209], stage057[234], stage056[241], stage055[258]}
   );
   gpc606_5 gpc606_5_6721(
      {stage055[211], stage055[212], stage055[213], stage055[214], stage055[215], stage055[216]},
      {stage057[190], stage057[191], stage057[192], stage057[193], stage057[194], stage057[195]},
      {stage059[268], stage058[210], stage057[235], stage056[242], stage055[259]}
   );
   gpc606_5 gpc606_5_6722(
      {stage055[217], stage055[218], stage055[219], stage055[220], stage055[221], stage055[222]},
      {stage057[196], stage057[197], stage057[198], stage057[199], stage057[200], stage057[201]},
      {stage059[269], stage058[211], stage057[236], stage056[243], stage055[260]}
   );
   gpc606_5 gpc606_5_6723(
      {stage055[223], stage055[224], stage055[225], stage055[226], stage055[227], stage055[228]},
      {stage057[202], stage057[203], stage057[204], stage057[205], stage057[206], stage057[207]},
      {stage059[270], stage058[212], stage057[237], stage056[244], stage055[261]}
   );
   gpc606_5 gpc606_5_6724(
      {stage055[229], stage055[230], stage055[231], stage055[232], stage055[233], stage055[234]},
      {stage057[208], stage057[209], stage057[210], stage057[211], stage057[212], stage057[213]},
      {stage059[271], stage058[213], stage057[238], stage056[245], stage055[262]}
   );
   gpc606_5 gpc606_5_6725(
      {stage055[235], stage055[236], stage055[237], stage055[238], stage055[239], stage055[240]},
      {stage057[214], stage057[215], stage057[216], stage057[217], stage057[218], stage057[219]},
      {stage059[272], stage058[214], stage057[239], stage056[246], stage055[263]}
   );
   gpc606_5 gpc606_5_6726(
      {stage055[241], stage055[242], stage055[243], stage055[244], stage055[245], stage055[246]},
      {stage057[220], stage057[221], stage057[222], stage057[223], stage057[224], stage057[225]},
      {stage059[273], stage058[215], stage057[240], stage056[247], stage055[264]}
   );
   gpc1_1 gpc1_1_6727(
      {stage056[205]},
      {stage056[248]}
   );
   gpc1_1 gpc1_1_6728(
      {stage056[206]},
      {stage056[249]}
   );
   gpc1_1 gpc1_1_6729(
      {stage056[207]},
      {stage056[250]}
   );
   gpc1_1 gpc1_1_6730(
      {stage056[208]},
      {stage056[251]}
   );
   gpc1_1 gpc1_1_6731(
      {stage056[209]},
      {stage056[252]}
   );
   gpc1_1 gpc1_1_6732(
      {stage056[210]},
      {stage056[253]}
   );
   gpc1_1 gpc1_1_6733(
      {stage056[211]},
      {stage056[254]}
   );
   gpc1_1 gpc1_1_6734(
      {stage056[212]},
      {stage056[255]}
   );
   gpc1_1 gpc1_1_6735(
      {stage056[213]},
      {stage056[256]}
   );
   gpc1_1 gpc1_1_6736(
      {stage056[214]},
      {stage056[257]}
   );
   gpc1_1 gpc1_1_6737(
      {stage056[215]},
      {stage056[258]}
   );
   gpc1_1 gpc1_1_6738(
      {stage056[216]},
      {stage056[259]}
   );
   gpc606_5 gpc606_5_6739(
      {stage056[217], stage056[218], stage056[219], stage056[220], stage056[221], stage056[222]},
      {stage058[180], stage058[181], stage058[182], stage058[183], stage058[184], stage058[185]},
      {stage060[215], stage059[274], stage058[216], stage057[241], stage056[260]}
   );
   gpc606_5 gpc606_5_6740(
      {stage056[223], stage056[224], stage056[225], stage056[226], stage056[227], stage056[228]},
      {stage058[186], stage058[187], stage058[188], stage058[189], stage058[190], stage058[191]},
      {stage060[216], stage059[275], stage058[217], stage057[242], stage056[261]}
   );
   gpc606_5 gpc606_5_6741(
      {stage056[229], stage056[230], stage056[231], stage056[232], stage056[233], stage056[234]},
      {stage058[192], stage058[193], stage058[194], stage058[195], stage058[196], stage058[197]},
      {stage060[217], stage059[276], stage058[218], stage057[243], stage056[262]}
   );
   gpc1_1 gpc1_1_6742(
      {stage057[226]},
      {stage057[244]}
   );
   gpc606_5 gpc606_5_6743(
      {stage057[227], stage057[228], stage057[229], stage057[230], stage057[231], stage057[232]},
      {stage059[216], stage059[217], stage059[218], stage059[219], stage059[220], stage059[221]},
      {stage061[246], stage060[218], stage059[277], stage058[219], stage057[245]}
   );
   gpc606_5 gpc606_5_6744(
      {stage058[198], stage058[199], stage058[200], stage058[201], stage058[202], stage058[203]},
      {stage060[190], stage060[191], stage060[192], stage060[193], stage060[194], stage060[195]},
      {stage062[215], stage061[247], stage060[219], stage059[278], stage058[220]}
   );
   gpc606_5 gpc606_5_6745(
      {stage058[204], stage058[205], stage058[206], stage058[207], stage058[208], 1'h0},
      {stage060[196], stage060[197], stage060[198], stage060[199], stage060[200], stage060[201]},
      {stage062[216], stage061[248], stage060[220], stage059[279], stage058[221]}
   );
   gpc1_1 gpc1_1_6746(
      {stage059[222]},
      {stage059[280]}
   );
   gpc1_1 gpc1_1_6747(
      {stage059[223]},
      {stage059[281]}
   );
   gpc1_1 gpc1_1_6748(
      {stage059[224]},
      {stage059[282]}
   );
   gpc1_1 gpc1_1_6749(
      {stage059[225]},
      {stage059[283]}
   );
   gpc1_1 gpc1_1_6750(
      {stage059[226]},
      {stage059[284]}
   );
   gpc1_1 gpc1_1_6751(
      {stage059[227]},
      {stage059[285]}
   );
   gpc1_1 gpc1_1_6752(
      {stage059[228]},
      {stage059[286]}
   );
   gpc1_1 gpc1_1_6753(
      {stage059[229]},
      {stage059[287]}
   );
   gpc1_1 gpc1_1_6754(
      {stage059[230]},
      {stage059[288]}
   );
   gpc1_1 gpc1_1_6755(
      {stage059[231]},
      {stage059[289]}
   );
   gpc615_5 gpc615_5_6756(
      {stage059[232], stage059[233], stage059[234], stage059[235], stage059[236]},
      {stage060[202]},
      {stage061[189], stage061[190], stage061[191], stage061[192], stage061[193], stage061[194]},
      {stage063[193], stage062[217], stage061[249], stage060[221], stage059[290]}
   );
   gpc615_5 gpc615_5_6757(
      {stage059[237], stage059[238], stage059[239], stage059[240], stage059[241]},
      {stage060[203]},
      {stage061[195], stage061[196], stage061[197], stage061[198], stage061[199], stage061[200]},
      {stage063[194], stage062[218], stage061[250], stage060[222], stage059[291]}
   );
   gpc615_5 gpc615_5_6758(
      {stage059[242], stage059[243], stage059[244], stage059[245], stage059[246]},
      {stage060[204]},
      {stage061[201], stage061[202], stage061[203], stage061[204], stage061[205], stage061[206]},
      {stage063[195], stage062[219], stage061[251], stage060[223], stage059[292]}
   );
   gpc615_5 gpc615_5_6759(
      {stage059[247], stage059[248], stage059[249], stage059[250], stage059[251]},
      {stage060[205]},
      {stage061[207], stage061[208], stage061[209], stage061[210], stage061[211], stage061[212]},
      {stage063[196], stage062[220], stage061[252], stage060[224], stage059[293]}
   );
   gpc615_5 gpc615_5_6760(
      {stage059[252], stage059[253], stage059[254], stage059[255], stage059[256]},
      {stage060[206]},
      {stage061[213], stage061[214], stage061[215], stage061[216], stage061[217], stage061[218]},
      {stage063[197], stage062[221], stage061[253], stage060[225], stage059[294]}
   );
   gpc615_5 gpc615_5_6761(
      {stage059[257], stage059[258], stage059[259], stage059[260], stage059[261]},
      {stage060[207]},
      {stage061[219], stage061[220], stage061[221], stage061[222], stage061[223], stage061[224]},
      {stage063[198], stage062[222], stage061[254], stage060[226], stage059[295]}
   );
   gpc615_5 gpc615_5_6762(
      {stage059[262], stage059[263], stage059[264], stage059[265], stage059[266]},
      {stage060[208]},
      {stage061[225], stage061[226], stage061[227], stage061[228], stage061[229], stage061[230]},
      {stage063[199], stage062[223], stage061[255], stage060[227], stage059[296]}
   );
   gpc606_5 gpc606_5_6763(
      {stage060[209], stage060[210], stage060[211], stage060[212], stage060[213], stage060[214]},
      {stage062[189], stage062[190], stage062[191], stage062[192], stage062[193], stage062[194]},
      {stage064[244], stage063[200], stage062[224], stage061[256], stage060[228]}
   );
   gpc1_1 gpc1_1_6764(
      {stage061[231]},
      {stage061[257]}
   );
   gpc1_1 gpc1_1_6765(
      {stage061[232]},
      {stage061[258]}
   );
   gpc1_1 gpc1_1_6766(
      {stage061[233]},
      {stage061[259]}
   );
   gpc606_5 gpc606_5_6767(
      {stage061[234], stage061[235], stage061[236], stage061[237], stage061[238], stage061[239]},
      {stage063[175], stage063[176], stage063[177], stage063[178], stage063[179], stage063[180]},
      {stage065[237], stage064[245], stage063[201], stage062[225], stage061[260]}
   );
   gpc606_5 gpc606_5_6768(
      {stage061[240], stage061[241], stage061[242], stage061[243], stage061[244], stage061[245]},
      {stage063[181], stage063[182], stage063[183], stage063[184], stage063[185], stage063[186]},
      {stage065[238], stage064[246], stage063[202], stage062[226], stage061[261]}
   );
   gpc1_1 gpc1_1_6769(
      {stage062[195]},
      {stage062[227]}
   );
   gpc1_1 gpc1_1_6770(
      {stage062[196]},
      {stage062[228]}
   );
   gpc1_1 gpc1_1_6771(
      {stage062[197]},
      {stage062[229]}
   );
   gpc1_1 gpc1_1_6772(
      {stage062[198]},
      {stage062[230]}
   );
   gpc1_1 gpc1_1_6773(
      {stage062[199]},
      {stage062[231]}
   );
   gpc1_1 gpc1_1_6774(
      {stage062[200]},
      {stage062[232]}
   );
   gpc1_1 gpc1_1_6775(
      {stage062[201]},
      {stage062[233]}
   );
   gpc1_1 gpc1_1_6776(
      {stage062[202]},
      {stage062[234]}
   );
   gpc1_1 gpc1_1_6777(
      {stage062[203]},
      {stage062[235]}
   );
   gpc1_1 gpc1_1_6778(
      {stage062[204]},
      {stage062[236]}
   );
   gpc615_5 gpc615_5_6779(
      {stage062[205], stage062[206], stage062[207], stage062[208], stage062[209]},
      {stage063[187]},
      {stage064[211], stage064[212], stage064[213], stage064[214], stage064[215], stage064[216]},
      {stage066[246], stage065[239], stage064[247], stage063[203], stage062[237]}
   );
   gpc615_5 gpc615_5_6780(
      {stage062[210], stage062[211], stage062[212], stage062[213], stage062[214]},
      {stage063[188]},
      {stage064[217], stage064[218], stage064[219], stage064[220], stage064[221], stage064[222]},
      {stage066[247], stage065[240], stage064[248], stage063[204], stage062[238]}
   );
   gpc1_1 gpc1_1_6781(
      {stage063[189]},
      {stage063[205]}
   );
   gpc1_1 gpc1_1_6782(
      {stage063[190]},
      {stage063[206]}
   );
   gpc1_1 gpc1_1_6783(
      {stage063[191]},
      {stage063[207]}
   );
   gpc1_1 gpc1_1_6784(
      {stage063[192]},
      {stage063[208]}
   );
   gpc1_1 gpc1_1_6785(
      {stage064[223]},
      {stage064[249]}
   );
   gpc1_1 gpc1_1_6786(
      {stage064[224]},
      {stage064[250]}
   );
   gpc1_1 gpc1_1_6787(
      {stage064[225]},
      {stage064[251]}
   );
   gpc1_1 gpc1_1_6788(
      {stage064[226]},
      {stage064[252]}
   );
   gpc1_1 gpc1_1_6789(
      {stage064[227]},
      {stage064[253]}
   );
   gpc606_5 gpc606_5_6790(
      {stage064[228], stage064[229], stage064[230], stage064[231], stage064[232], stage064[233]},
      {stage066[211], stage066[212], stage066[213], stage066[214], stage066[215], stage066[216]},
      {stage068[241], stage067[244], stage066[248], stage065[241], stage064[254]}
   );
   gpc615_5 gpc615_5_6791(
      {stage064[234], stage064[235], stage064[236], stage064[237], stage064[238]},
      {stage065[199]},
      {stage066[217], stage066[218], stage066[219], stage066[220], stage066[221], stage066[222]},
      {stage068[242], stage067[245], stage066[249], stage065[242], stage064[255]}
   );
   gpc615_5 gpc615_5_6792(
      {stage064[239], stage064[240], stage064[241], stage064[242], stage064[243]},
      {stage065[200]},
      {stage066[223], stage066[224], stage066[225], stage066[226], stage066[227], stage066[228]},
      {stage068[243], stage067[246], stage066[250], stage065[243], stage064[256]}
   );
   gpc1_1 gpc1_1_6793(
      {stage065[201]},
      {stage065[244]}
   );
   gpc1_1 gpc1_1_6794(
      {stage065[202]},
      {stage065[245]}
   );
   gpc1_1 gpc1_1_6795(
      {stage065[203]},
      {stage065[246]}
   );
   gpc1_1 gpc1_1_6796(
      {stage065[204]},
      {stage065[247]}
   );
   gpc1_1 gpc1_1_6797(
      {stage065[205]},
      {stage065[248]}
   );
   gpc1_1 gpc1_1_6798(
      {stage065[206]},
      {stage065[249]}
   );
   gpc606_5 gpc606_5_6799(
      {stage065[207], stage065[208], stage065[209], stage065[210], stage065[211], stage065[212]},
      {stage067[213], stage067[214], stage067[215], stage067[216], stage067[217], stage067[218]},
      {stage069[233], stage068[244], stage067[247], stage066[251], stage065[250]}
   );
   gpc606_5 gpc606_5_6800(
      {stage065[213], stage065[214], stage065[215], stage065[216], stage065[217], stage065[218]},
      {stage067[219], stage067[220], stage067[221], stage067[222], stage067[223], stage067[224]},
      {stage069[234], stage068[245], stage067[248], stage066[252], stage065[251]}
   );
   gpc606_5 gpc606_5_6801(
      {stage065[219], stage065[220], stage065[221], stage065[222], stage065[223], stage065[224]},
      {stage067[225], stage067[226], stage067[227], stage067[228], stage067[229], stage067[230]},
      {stage069[235], stage068[246], stage067[249], stage066[253], stage065[252]}
   );
   gpc606_5 gpc606_5_6802(
      {stage065[225], stage065[226], stage065[227], stage065[228], stage065[229], stage065[230]},
      {stage067[231], stage067[232], stage067[233], stage067[234], stage067[235], stage067[236]},
      {stage069[236], stage068[247], stage067[250], stage066[254], stage065[253]}
   );
   gpc606_5 gpc606_5_6803(
      {stage065[231], stage065[232], stage065[233], stage065[234], stage065[235], stage065[236]},
      {stage067[237], stage067[238], stage067[239], stage067[240], stage067[241], stage067[242]},
      {stage069[237], stage068[248], stage067[251], stage066[255], stage065[254]}
   );
   gpc1_1 gpc1_1_6804(
      {stage066[229]},
      {stage066[256]}
   );
   gpc1_1 gpc1_1_6805(
      {stage066[230]},
      {stage066[257]}
   );
   gpc1_1 gpc1_1_6806(
      {stage066[231]},
      {stage066[258]}
   );
   gpc1_1 gpc1_1_6807(
      {stage066[232]},
      {stage066[259]}
   );
   gpc1_1 gpc1_1_6808(
      {stage066[233]},
      {stage066[260]}
   );
   gpc1_1 gpc1_1_6809(
      {stage066[234]},
      {stage066[261]}
   );
   gpc1_1 gpc1_1_6810(
      {stage066[235]},
      {stage066[262]}
   );
   gpc1_1 gpc1_1_6811(
      {stage066[236]},
      {stage066[263]}
   );
   gpc1_1 gpc1_1_6812(
      {stage066[237]},
      {stage066[264]}
   );
   gpc1_1 gpc1_1_6813(
      {stage066[238]},
      {stage066[265]}
   );
   gpc1_1 gpc1_1_6814(
      {stage066[239]},
      {stage066[266]}
   );
   gpc1_1 gpc1_1_6815(
      {stage066[240]},
      {stage066[267]}
   );
   gpc1_1 gpc1_1_6816(
      {stage066[241]},
      {stage066[268]}
   );
   gpc1_1 gpc1_1_6817(
      {stage066[242]},
      {stage066[269]}
   );
   gpc1_1 gpc1_1_6818(
      {stage066[243]},
      {stage066[270]}
   );
   gpc1_1 gpc1_1_6819(
      {stage066[244]},
      {stage066[271]}
   );
   gpc1_1 gpc1_1_6820(
      {stage066[245]},
      {stage066[272]}
   );
   gpc1_1 gpc1_1_6821(
      {stage067[243]},
      {stage067[252]}
   );
   gpc1_1 gpc1_1_6822(
      {stage068[210]},
      {stage068[249]}
   );
   gpc1_1 gpc1_1_6823(
      {stage068[211]},
      {stage068[250]}
   );
   gpc1_1 gpc1_1_6824(
      {stage068[212]},
      {stage068[251]}
   );
   gpc1_1 gpc1_1_6825(
      {stage068[213]},
      {stage068[252]}
   );
   gpc1_1 gpc1_1_6826(
      {stage068[214]},
      {stage068[253]}
   );
   gpc1_1 gpc1_1_6827(
      {stage068[215]},
      {stage068[254]}
   );
   gpc1_1 gpc1_1_6828(
      {stage068[216]},
      {stage068[255]}
   );
   gpc1_1 gpc1_1_6829(
      {stage068[217]},
      {stage068[256]}
   );
   gpc1_1 gpc1_1_6830(
      {stage068[218]},
      {stage068[257]}
   );
   gpc1_1 gpc1_1_6831(
      {stage068[219]},
      {stage068[258]}
   );
   gpc623_5 gpc623_5_6832(
      {stage068[220], stage068[221], stage068[222]},
      {stage069[183], stage069[184]},
      {stage070[189], stage070[190], stage070[191], stage070[192], stage070[193], stage070[194]},
      {stage072[267], stage071[237], stage070[234], stage069[238], stage068[259]}
   );
   gpc623_5 gpc623_5_6833(
      {stage068[223], stage068[224], stage068[225]},
      {stage069[185], stage069[186]},
      {stage070[195], stage070[196], stage070[197], stage070[198], stage070[199], stage070[200]},
      {stage072[268], stage071[238], stage070[235], stage069[239], stage068[260]}
   );
   gpc623_5 gpc623_5_6834(
      {stage068[226], stage068[227], stage068[228]},
      {stage069[187], stage069[188]},
      {stage070[201], stage070[202], stage070[203], stage070[204], stage070[205], stage070[206]},
      {stage072[269], stage071[239], stage070[236], stage069[240], stage068[261]}
   );
   gpc623_5 gpc623_5_6835(
      {stage068[229], stage068[230], stage068[231]},
      {stage069[189], stage069[190]},
      {stage070[207], stage070[208], stage070[209], stage070[210], stage070[211], stage070[212]},
      {stage072[270], stage071[240], stage070[237], stage069[241], stage068[262]}
   );
   gpc623_5 gpc623_5_6836(
      {stage068[232], stage068[233], stage068[234]},
      {stage069[191], stage069[192]},
      {stage070[213], stage070[214], stage070[215], stage070[216], stage070[217], stage070[218]},
      {stage072[271], stage071[241], stage070[238], stage069[242], stage068[263]}
   );
   gpc623_5 gpc623_5_6837(
      {stage068[235], stage068[236], stage068[237]},
      {stage069[193], stage069[194]},
      {stage070[219], stage070[220], stage070[221], stage070[222], stage070[223], stage070[224]},
      {stage072[272], stage071[242], stage070[239], stage069[243], stage068[264]}
   );
   gpc623_5 gpc623_5_6838(
      {stage068[238], stage068[239], stage068[240]},
      {stage069[195], stage069[196]},
      {stage070[225], stage070[226], stage070[227], stage070[228], stage070[229], stage070[230]},
      {stage072[273], stage071[243], stage070[240], stage069[244], stage068[265]}
   );
   gpc1_1 gpc1_1_6839(
      {stage069[197]},
      {stage069[245]}
   );
   gpc1_1 gpc1_1_6840(
      {stage069[198]},
      {stage069[246]}
   );
   gpc1_1 gpc1_1_6841(
      {stage069[199]},
      {stage069[247]}
   );
   gpc1_1 gpc1_1_6842(
      {stage069[200]},
      {stage069[248]}
   );
   gpc1_1 gpc1_1_6843(
      {stage069[201]},
      {stage069[249]}
   );
   gpc1_1 gpc1_1_6844(
      {stage069[202]},
      {stage069[250]}
   );
   gpc606_5 gpc606_5_6845(
      {stage069[203], stage069[204], stage069[205], stage069[206], stage069[207], stage069[208]},
      {stage071[188], stage071[189], stage071[190], stage071[191], stage071[192], stage071[193]},
      {stage073[217], stage072[274], stage071[244], stage070[241], stage069[251]}
   );
   gpc606_5 gpc606_5_6846(
      {stage069[209], stage069[210], stage069[211], stage069[212], stage069[213], stage069[214]},
      {stage071[194], stage071[195], stage071[196], stage071[197], stage071[198], stage071[199]},
      {stage073[218], stage072[275], stage071[245], stage070[242], stage069[252]}
   );
   gpc606_5 gpc606_5_6847(
      {stage069[215], stage069[216], stage069[217], stage069[218], stage069[219], stage069[220]},
      {stage071[200], stage071[201], stage071[202], stage071[203], stage071[204], stage071[205]},
      {stage073[219], stage072[276], stage071[246], stage070[243], stage069[253]}
   );
   gpc606_5 gpc606_5_6848(
      {stage069[221], stage069[222], stage069[223], stage069[224], stage069[225], stage069[226]},
      {stage071[206], stage071[207], stage071[208], stage071[209], stage071[210], stage071[211]},
      {stage073[220], stage072[277], stage071[247], stage070[244], stage069[254]}
   );
   gpc606_5 gpc606_5_6849(
      {stage069[227], stage069[228], stage069[229], stage069[230], stage069[231], stage069[232]},
      {stage071[212], stage071[213], stage071[214], stage071[215], stage071[216], stage071[217]},
      {stage073[221], stage072[278], stage071[248], stage070[245], stage069[255]}
   );
   gpc1_1 gpc1_1_6850(
      {stage070[231]},
      {stage070[246]}
   );
   gpc1_1 gpc1_1_6851(
      {stage070[232]},
      {stage070[247]}
   );
   gpc1_1 gpc1_1_6852(
      {stage070[233]},
      {stage070[248]}
   );
   gpc1_1 gpc1_1_6853(
      {stage071[218]},
      {stage071[249]}
   );
   gpc1_1 gpc1_1_6854(
      {stage071[219]},
      {stage071[250]}
   );
   gpc1_1 gpc1_1_6855(
      {stage071[220]},
      {stage071[251]}
   );
   gpc1_1 gpc1_1_6856(
      {stage071[221]},
      {stage071[252]}
   );
   gpc615_5 gpc615_5_6857(
      {stage071[222], stage071[223], stage071[224], stage071[225], stage071[226]},
      {stage072[222]},
      {stage073[193], stage073[194], stage073[195], stage073[196], stage073[197], stage073[198]},
      {stage075[193], stage074[227], stage073[222], stage072[279], stage071[253]}
   );
   gpc615_5 gpc615_5_6858(
      {stage071[227], stage071[228], stage071[229], stage071[230], stage071[231]},
      {stage072[223]},
      {stage073[199], stage073[200], stage073[201], stage073[202], stage073[203], stage073[204]},
      {stage075[194], stage074[228], stage073[223], stage072[280], stage071[254]}
   );
   gpc615_5 gpc615_5_6859(
      {stage071[232], stage071[233], stage071[234], stage071[235], stage071[236]},
      {stage072[224]},
      {stage073[205], stage073[206], stage073[207], stage073[208], stage073[209], stage073[210]},
      {stage075[195], stage074[229], stage073[224], stage072[281], stage071[255]}
   );
   gpc1_1 gpc1_1_6860(
      {stage072[225]},
      {stage072[282]}
   );
   gpc1_1 gpc1_1_6861(
      {stage072[226]},
      {stage072[283]}
   );
   gpc1_1 gpc1_1_6862(
      {stage072[227]},
      {stage072[284]}
   );
   gpc1_1 gpc1_1_6863(
      {stage072[228]},
      {stage072[285]}
   );
   gpc1_1 gpc1_1_6864(
      {stage072[229]},
      {stage072[286]}
   );
   gpc1_1 gpc1_1_6865(
      {stage072[230]},
      {stage072[287]}
   );
   gpc1_1 gpc1_1_6866(
      {stage072[231]},
      {stage072[288]}
   );
   gpc1_1 gpc1_1_6867(
      {stage072[232]},
      {stage072[289]}
   );
   gpc1_1 gpc1_1_6868(
      {stage072[233]},
      {stage072[290]}
   );
   gpc1_1 gpc1_1_6869(
      {stage072[234]},
      {stage072[291]}
   );
   gpc1_1 gpc1_1_6870(
      {stage072[235]},
      {stage072[292]}
   );
   gpc1_1 gpc1_1_6871(
      {stage072[236]},
      {stage072[293]}
   );
   gpc606_5 gpc606_5_6872(
      {stage072[237], stage072[238], stage072[239], stage072[240], stage072[241], stage072[242]},
      {stage074[189], stage074[190], stage074[191], stage074[192], stage074[193], stage074[194]},
      {stage076[197], stage075[196], stage074[230], stage073[225], stage072[294]}
   );
   gpc606_5 gpc606_5_6873(
      {stage072[243], stage072[244], stage072[245], stage072[246], stage072[247], stage072[248]},
      {stage074[195], stage074[196], stage074[197], stage074[198], stage074[199], stage074[200]},
      {stage076[198], stage075[197], stage074[231], stage073[226], stage072[295]}
   );
   gpc606_5 gpc606_5_6874(
      {stage072[249], stage072[250], stage072[251], stage072[252], stage072[253], stage072[254]},
      {stage074[201], stage074[202], stage074[203], stage074[204], stage074[205], stage074[206]},
      {stage076[199], stage075[198], stage074[232], stage073[227], stage072[296]}
   );
   gpc606_5 gpc606_5_6875(
      {stage072[255], stage072[256], stage072[257], stage072[258], stage072[259], stage072[260]},
      {stage074[207], stage074[208], stage074[209], stage074[210], stage074[211], stage074[212]},
      {stage076[200], stage075[199], stage074[233], stage073[228], stage072[297]}
   );
   gpc606_5 gpc606_5_6876(
      {stage072[261], stage072[262], stage072[263], stage072[264], stage072[265], stage072[266]},
      {stage074[213], stage074[214], stage074[215], stage074[216], stage074[217], stage074[218]},
      {stage076[201], stage075[200], stage074[234], stage073[229], stage072[298]}
   );
   gpc1_1 gpc1_1_6877(
      {stage073[211]},
      {stage073[230]}
   );
   gpc615_5 gpc615_5_6878(
      {stage073[212], stage073[213], stage073[214], stage073[215], stage073[216]},
      {stage074[219]},
      {stage075[169], stage075[170], stage075[171], stage075[172], stage075[173], stage075[174]},
      {stage077[230], stage076[202], stage075[201], stage074[235], stage073[231]}
   );
   gpc1_1 gpc1_1_6879(
      {stage074[220]},
      {stage074[236]}
   );
   gpc1_1 gpc1_1_6880(
      {stage074[221]},
      {stage074[237]}
   );
   gpc1_1 gpc1_1_6881(
      {stage074[222]},
      {stage074[238]}
   );
   gpc1_1 gpc1_1_6882(
      {stage074[223]},
      {stage074[239]}
   );
   gpc1_1 gpc1_1_6883(
      {stage074[224]},
      {stage074[240]}
   );
   gpc1_1 gpc1_1_6884(
      {stage074[225]},
      {stage074[241]}
   );
   gpc1_1 gpc1_1_6885(
      {stage074[226]},
      {stage074[242]}
   );
   gpc606_5 gpc606_5_6886(
      {stage075[175], stage075[176], stage075[177], stage075[178], stage075[179], stage075[180]},
      {stage077[203], stage077[204], stage077[205], stage077[206], stage077[207], stage077[208]},
      {stage079[216], stage078[207], stage077[231], stage076[203], stage075[202]}
   );
   gpc606_5 gpc606_5_6887(
      {stage075[181], stage075[182], stage075[183], stage075[184], stage075[185], stage075[186]},
      {stage077[209], stage077[210], stage077[211], stage077[212], stage077[213], stage077[214]},
      {stage079[217], stage078[208], stage077[232], stage076[204], stage075[203]}
   );
   gpc606_5 gpc606_5_6888(
      {stage075[187], stage075[188], stage075[189], stage075[190], stage075[191], stage075[192]},
      {stage077[215], stage077[216], stage077[217], stage077[218], stage077[219], stage077[220]},
      {stage079[218], stage078[209], stage077[233], stage076[205], stage075[204]}
   );
   gpc615_5 gpc615_5_6889(
      {stage076[182], stage076[183], stage076[184], stage076[185], stage076[186]},
      {stage077[221]},
      {stage078[174], stage078[175], stage078[176], stage078[177], stage078[178], stage078[179]},
      {stage080[232], stage079[219], stage078[210], stage077[234], stage076[206]}
   );
   gpc615_5 gpc615_5_6890(
      {stage076[187], stage076[188], stage076[189], stage076[190], stage076[191]},
      {stage077[222]},
      {stage078[180], stage078[181], stage078[182], stage078[183], stage078[184], stage078[185]},
      {stage080[233], stage079[220], stage078[211], stage077[235], stage076[207]}
   );
   gpc615_5 gpc615_5_6891(
      {stage076[192], stage076[193], stage076[194], stage076[195], stage076[196]},
      {stage077[223]},
      {stage078[186], stage078[187], stage078[188], stage078[189], stage078[190], stage078[191]},
      {stage080[234], stage079[221], stage078[212], stage077[236], stage076[208]}
   );
   gpc1_1 gpc1_1_6892(
      {stage077[224]},
      {stage077[237]}
   );
   gpc1_1 gpc1_1_6893(
      {stage077[225]},
      {stage077[238]}
   );
   gpc1_1 gpc1_1_6894(
      {stage077[226]},
      {stage077[239]}
   );
   gpc1_1 gpc1_1_6895(
      {stage077[227]},
      {stage077[240]}
   );
   gpc1_1 gpc1_1_6896(
      {stage077[228]},
      {stage077[241]}
   );
   gpc1_1 gpc1_1_6897(
      {stage077[229]},
      {stage077[242]}
   );
   gpc1_1 gpc1_1_6898(
      {stage078[192]},
      {stage078[213]}
   );
   gpc1_1 gpc1_1_6899(
      {stage078[193]},
      {stage078[214]}
   );
   gpc1_1 gpc1_1_6900(
      {stage078[194]},
      {stage078[215]}
   );
   gpc1_1 gpc1_1_6901(
      {stage078[195]},
      {stage078[216]}
   );
   gpc1_1 gpc1_1_6902(
      {stage078[196]},
      {stage078[217]}
   );
   gpc1_1 gpc1_1_6903(
      {stage078[197]},
      {stage078[218]}
   );
   gpc1_1 gpc1_1_6904(
      {stage078[198]},
      {stage078[219]}
   );
   gpc1_1 gpc1_1_6905(
      {stage078[199]},
      {stage078[220]}
   );
   gpc1_1 gpc1_1_6906(
      {stage078[200]},
      {stage078[221]}
   );
   gpc1_1 gpc1_1_6907(
      {stage078[201]},
      {stage078[222]}
   );
   gpc1_1 gpc1_1_6908(
      {stage078[202]},
      {stage078[223]}
   );
   gpc1_1 gpc1_1_6909(
      {stage078[203]},
      {stage078[224]}
   );
   gpc1_1 gpc1_1_6910(
      {stage078[204]},
      {stage078[225]}
   );
   gpc1_1 gpc1_1_6911(
      {stage078[205]},
      {stage078[226]}
   );
   gpc1_1 gpc1_1_6912(
      {stage078[206]},
      {stage078[227]}
   );
   gpc1_1 gpc1_1_6913(
      {stage079[187]},
      {stage079[222]}
   );
   gpc1_1 gpc1_1_6914(
      {stage079[188]},
      {stage079[223]}
   );
   gpc1_1 gpc1_1_6915(
      {stage079[189]},
      {stage079[224]}
   );
   gpc1_1 gpc1_1_6916(
      {stage079[190]},
      {stage079[225]}
   );
   gpc1_1 gpc1_1_6917(
      {stage079[191]},
      {stage079[226]}
   );
   gpc1_1 gpc1_1_6918(
      {stage079[192]},
      {stage079[227]}
   );
   gpc1_1 gpc1_1_6919(
      {stage079[193]},
      {stage079[228]}
   );
   gpc1_1 gpc1_1_6920(
      {stage079[194]},
      {stage079[229]}
   );
   gpc1_1 gpc1_1_6921(
      {stage079[195]},
      {stage079[230]}
   );
   gpc1_1 gpc1_1_6922(
      {stage079[196]},
      {stage079[231]}
   );
   gpc1_1 gpc1_1_6923(
      {stage079[197]},
      {stage079[232]}
   );
   gpc1_1 gpc1_1_6924(
      {stage079[198]},
      {stage079[233]}
   );
   gpc1_1 gpc1_1_6925(
      {stage079[199]},
      {stage079[234]}
   );
   gpc606_5 gpc606_5_6926(
      {stage079[200], stage079[201], stage079[202], stage079[203], stage079[204], stage079[205]},
      {stage081[175], stage081[176], stage081[177], stage081[178], stage081[179], stage081[180]},
      {stage083[246], stage082[240], stage081[238], stage080[235], stage079[235]}
   );
   gpc615_5 gpc615_5_6927(
      {stage079[206], stage079[207], stage079[208], stage079[209], stage079[210]},
      {stage080[203]},
      {stage081[181], stage081[182], stage081[183], stage081[184], stage081[185], stage081[186]},
      {stage083[247], stage082[241], stage081[239], stage080[236], stage079[236]}
   );
   gpc615_5 gpc615_5_6928(
      {stage079[211], stage079[212], stage079[213], stage079[214], stage079[215]},
      {stage080[204]},
      {stage081[187], stage081[188], stage081[189], stage081[190], stage081[191], stage081[192]},
      {stage083[248], stage082[242], stage081[240], stage080[237], stage079[237]}
   );
   gpc1_1 gpc1_1_6929(
      {stage080[205]},
      {stage080[238]}
   );
   gpc1_1 gpc1_1_6930(
      {stage080[206]},
      {stage080[239]}
   );
   gpc1_1 gpc1_1_6931(
      {stage080[207]},
      {stage080[240]}
   );
   gpc1_1 gpc1_1_6932(
      {stage080[208]},
      {stage080[241]}
   );
   gpc1_1 gpc1_1_6933(
      {stage080[209]},
      {stage080[242]}
   );
   gpc1_1 gpc1_1_6934(
      {stage080[210]},
      {stage080[243]}
   );
   gpc1_1 gpc1_1_6935(
      {stage080[211]},
      {stage080[244]}
   );
   gpc1_1 gpc1_1_6936(
      {stage080[212]},
      {stage080[245]}
   );
   gpc1_1 gpc1_1_6937(
      {stage080[213]},
      {stage080[246]}
   );
   gpc1_1 gpc1_1_6938(
      {stage080[214]},
      {stage080[247]}
   );
   gpc1_1 gpc1_1_6939(
      {stage080[215]},
      {stage080[248]}
   );
   gpc1_1 gpc1_1_6940(
      {stage080[216]},
      {stage080[249]}
   );
   gpc615_5 gpc615_5_6941(
      {stage080[217], stage080[218], stage080[219], stage080[220], stage080[221]},
      {stage081[193]},
      {stage082[215], stage082[216], stage082[217], stage082[218], stage082[219], stage082[220]},
      {stage084[218], stage083[249], stage082[243], stage081[241], stage080[250]}
   );
   gpc615_5 gpc615_5_6942(
      {stage080[222], stage080[223], stage080[224], stage080[225], stage080[226]},
      {stage081[194]},
      {stage082[221], stage082[222], stage082[223], stage082[224], stage082[225], stage082[226]},
      {stage084[219], stage083[250], stage082[244], stage081[242], stage080[251]}
   );
   gpc615_5 gpc615_5_6943(
      {stage080[227], stage080[228], stage080[229], stage080[230], stage080[231]},
      {stage081[195]},
      {stage082[227], stage082[228], stage082[229], stage082[230], stage082[231], stage082[232]},
      {stage084[220], stage083[251], stage082[245], stage081[243], stage080[252]}
   );
   gpc1_1 gpc1_1_6944(
      {stage081[196]},
      {stage081[244]}
   );
   gpc1_1 gpc1_1_6945(
      {stage081[197]},
      {stage081[245]}
   );
   gpc1_1 gpc1_1_6946(
      {stage081[198]},
      {stage081[246]}
   );
   gpc1_1 gpc1_1_6947(
      {stage081[199]},
      {stage081[247]}
   );
   gpc1_1 gpc1_1_6948(
      {stage081[200]},
      {stage081[248]}
   );
   gpc1_1 gpc1_1_6949(
      {stage081[201]},
      {stage081[249]}
   );
   gpc1_1 gpc1_1_6950(
      {stage081[202]},
      {stage081[250]}
   );
   gpc1_1 gpc1_1_6951(
      {stage081[203]},
      {stage081[251]}
   );
   gpc606_5 gpc606_5_6952(
      {stage081[204], stage081[205], stage081[206], stage081[207], stage081[208], stage081[209]},
      {stage083[196], stage083[197], stage083[198], stage083[199], stage083[200], stage083[201]},
      {stage085[249], stage084[221], stage083[252], stage082[246], stage081[252]}
   );
   gpc606_5 gpc606_5_6953(
      {stage081[210], stage081[211], stage081[212], stage081[213], stage081[214], stage081[215]},
      {stage083[202], stage083[203], stage083[204], stage083[205], stage083[206], stage083[207]},
      {stage085[250], stage084[222], stage083[253], stage082[247], stage081[253]}
   );
   gpc606_5 gpc606_5_6954(
      {stage081[216], stage081[217], stage081[218], stage081[219], stage081[220], stage081[221]},
      {stage083[208], stage083[209], stage083[210], stage083[211], stage083[212], stage083[213]},
      {stage085[251], stage084[223], stage083[254], stage082[248], stage081[254]}
   );
   gpc606_5 gpc606_5_6955(
      {stage081[222], stage081[223], stage081[224], stage081[225], stage081[226], stage081[227]},
      {stage083[214], stage083[215], stage083[216], stage083[217], stage083[218], stage083[219]},
      {stage085[252], stage084[224], stage083[255], stage082[249], stage081[255]}
   );
   gpc615_5 gpc615_5_6956(
      {stage081[228], stage081[229], stage081[230], stage081[231], stage081[232]},
      {stage082[233]},
      {stage083[220], stage083[221], stage083[222], stage083[223], stage083[224], stage083[225]},
      {stage085[253], stage084[225], stage083[256], stage082[250], stage081[256]}
   );
   gpc615_5 gpc615_5_6957(
      {stage081[233], stage081[234], stage081[235], stage081[236], stage081[237]},
      {stage082[234]},
      {stage083[226], stage083[227], stage083[228], stage083[229], stage083[230], stage083[231]},
      {stage085[254], stage084[226], stage083[257], stage082[251], stage081[257]}
   );
   gpc1_1 gpc1_1_6958(
      {stage082[235]},
      {stage082[252]}
   );
   gpc1_1 gpc1_1_6959(
      {stage082[236]},
      {stage082[253]}
   );
   gpc623_5 gpc623_5_6960(
      {stage082[237], stage082[238], stage082[239]},
      {stage083[232], stage083[233]},
      {stage084[197], stage084[198], stage084[199], stage084[200], stage084[201], stage084[202]},
      {stage086[243], stage085[255], stage084[227], stage083[258], stage082[254]}
   );
   gpc606_5 gpc606_5_6961(
      {stage083[234], stage083[235], stage083[236], stage083[237], stage083[238], stage083[239]},
      {stage085[218], stage085[219], stage085[220], stage085[221], stage085[222], stage085[223]},
      {stage087[213], stage086[244], stage085[256], stage084[228], stage083[259]}
   );
   gpc606_5 gpc606_5_6962(
      {stage083[240], stage083[241], stage083[242], stage083[243], stage083[244], stage083[245]},
      {stage085[224], stage085[225], stage085[226], stage085[227], stage085[228], stage085[229]},
      {stage087[214], stage086[245], stage085[257], stage084[229], stage083[260]}
   );
   gpc1_1 gpc1_1_6963(
      {stage084[203]},
      {stage084[230]}
   );
   gpc1_1 gpc1_1_6964(
      {stage084[204]},
      {stage084[231]}
   );
   gpc1_1 gpc1_1_6965(
      {stage084[205]},
      {stage084[232]}
   );
   gpc606_5 gpc606_5_6966(
      {stage084[206], stage084[207], stage084[208], stage084[209], stage084[210], stage084[211]},
      {stage086[205], stage086[206], stage086[207], stage086[208], stage086[209], stage086[210]},
      {stage088[246], stage087[215], stage086[246], stage085[258], stage084[233]}
   );
   gpc606_5 gpc606_5_6967(
      {stage084[212], stage084[213], stage084[214], stage084[215], stage084[216], stage084[217]},
      {stage086[211], stage086[212], stage086[213], stage086[214], stage086[215], stage086[216]},
      {stage088[247], stage087[216], stage086[247], stage085[259], stage084[234]}
   );
   gpc1_1 gpc1_1_6968(
      {stage085[230]},
      {stage085[260]}
   );
   gpc1_1 gpc1_1_6969(
      {stage085[231]},
      {stage085[261]}
   );
   gpc606_5 gpc606_5_6970(
      {stage085[232], stage085[233], stage085[234], stage085[235], stage085[236], stage085[237]},
      {stage087[183], stage087[184], stage087[185], stage087[186], stage087[187], stage087[188]},
      {stage089[216], stage088[248], stage087[217], stage086[248], stage085[262]}
   );
   gpc606_5 gpc606_5_6971(
      {stage085[238], stage085[239], stage085[240], stage085[241], stage085[242], stage085[243]},
      {stage087[189], stage087[190], stage087[191], stage087[192], stage087[193], stage087[194]},
      {stage089[217], stage088[249], stage087[218], stage086[249], stage085[263]}
   );
   gpc615_5 gpc615_5_6972(
      {stage085[244], stage085[245], stage085[246], stage085[247], stage085[248]},
      {stage086[217]},
      {stage087[195], stage087[196], stage087[197], stage087[198], stage087[199], stage087[200]},
      {stage089[218], stage088[250], stage087[219], stage086[250], stage085[264]}
   );
   gpc1_1 gpc1_1_6973(
      {stage086[218]},
      {stage086[251]}
   );
   gpc1_1 gpc1_1_6974(
      {stage086[219]},
      {stage086[252]}
   );
   gpc1_1 gpc1_1_6975(
      {stage086[220]},
      {stage086[253]}
   );
   gpc1_1 gpc1_1_6976(
      {stage086[221]},
      {stage086[254]}
   );
   gpc1_1 gpc1_1_6977(
      {stage086[222]},
      {stage086[255]}
   );
   gpc1_1 gpc1_1_6978(
      {stage086[223]},
      {stage086[256]}
   );
   gpc1_1 gpc1_1_6979(
      {stage086[224]},
      {stage086[257]}
   );
   gpc1_1 gpc1_1_6980(
      {stage086[225]},
      {stage086[258]}
   );
   gpc1_1 gpc1_1_6981(
      {stage086[226]},
      {stage086[259]}
   );
   gpc1_1 gpc1_1_6982(
      {stage086[227]},
      {stage086[260]}
   );
   gpc1_1 gpc1_1_6983(
      {stage086[228]},
      {stage086[261]}
   );
   gpc1_1 gpc1_1_6984(
      {stage086[229]},
      {stage086[262]}
   );
   gpc1_1 gpc1_1_6985(
      {stage086[230]},
      {stage086[263]}
   );
   gpc1_1 gpc1_1_6986(
      {stage086[231]},
      {stage086[264]}
   );
   gpc1_1 gpc1_1_6987(
      {stage086[232]},
      {stage086[265]}
   );
   gpc1_1 gpc1_1_6988(
      {stage086[233]},
      {stage086[266]}
   );
   gpc1_1 gpc1_1_6989(
      {stage086[234]},
      {stage086[267]}
   );
   gpc1_1 gpc1_1_6990(
      {stage086[235]},
      {stage086[268]}
   );
   gpc1_1 gpc1_1_6991(
      {stage086[236]},
      {stage086[269]}
   );
   gpc606_5 gpc606_5_6992(
      {stage086[237], stage086[238], stage086[239], stage086[240], stage086[241], stage086[242]},
      {stage088[220], stage088[221], stage088[222], stage088[223], stage088[224], stage088[225]},
      {stage090[217], stage089[219], stage088[251], stage087[220], stage086[270]}
   );
   gpc606_5 gpc606_5_6993(
      {stage087[201], stage087[202], stage087[203], stage087[204], stage087[205], stage087[206]},
      {stage089[166], stage089[167], stage089[168], stage089[169], stage089[170], stage089[171]},
      {stage091[255], stage090[218], stage089[220], stage088[252], stage087[221]}
   );
   gpc606_5 gpc606_5_6994(
      {stage087[207], stage087[208], stage087[209], stage087[210], stage087[211], stage087[212]},
      {stage089[172], stage089[173], stage089[174], stage089[175], stage089[176], stage089[177]},
      {stage091[256], stage090[219], stage089[221], stage088[253], stage087[222]}
   );
   gpc1_1 gpc1_1_6995(
      {stage088[226]},
      {stage088[254]}
   );
   gpc1_1 gpc1_1_6996(
      {stage088[227]},
      {stage088[255]}
   );
   gpc1_1 gpc1_1_6997(
      {stage088[228]},
      {stage088[256]}
   );
   gpc1_1 gpc1_1_6998(
      {stage088[229]},
      {stage088[257]}
   );
   gpc1_1 gpc1_1_6999(
      {stage088[230]},
      {stage088[258]}
   );
   gpc1_1 gpc1_1_7000(
      {stage088[231]},
      {stage088[259]}
   );
   gpc1_1 gpc1_1_7001(
      {stage088[232]},
      {stage088[260]}
   );
   gpc1_1 gpc1_1_7002(
      {stage088[233]},
      {stage088[261]}
   );
   gpc606_5 gpc606_5_7003(
      {stage088[234], stage088[235], stage088[236], stage088[237], stage088[238], stage088[239]},
      {stage090[180], stage090[181], stage090[182], stage090[183], stage090[184], stage090[185]},
      {stage092[227], stage091[257], stage090[220], stage089[222], stage088[262]}
   );
   gpc606_5 gpc606_5_7004(
      {stage088[240], stage088[241], stage088[242], stage088[243], stage088[244], stage088[245]},
      {stage090[186], stage090[187], stage090[188], stage090[189], stage090[190], stage090[191]},
      {stage092[228], stage091[258], stage090[221], stage089[223], stage088[263]}
   );
   gpc1_1 gpc1_1_7005(
      {stage089[178]},
      {stage089[224]}
   );
   gpc1_1 gpc1_1_7006(
      {stage089[179]},
      {stage089[225]}
   );
   gpc1_1 gpc1_1_7007(
      {stage089[180]},
      {stage089[226]}
   );
   gpc1_1 gpc1_1_7008(
      {stage089[181]},
      {stage089[227]}
   );
   gpc1_1 gpc1_1_7009(
      {stage089[182]},
      {stage089[228]}
   );
   gpc1_1 gpc1_1_7010(
      {stage089[183]},
      {stage089[229]}
   );
   gpc1_1 gpc1_1_7011(
      {stage089[184]},
      {stage089[230]}
   );
   gpc1_1 gpc1_1_7012(
      {stage089[185]},
      {stage089[231]}
   );
   gpc1_1 gpc1_1_7013(
      {stage089[186]},
      {stage089[232]}
   );
   gpc1_1 gpc1_1_7014(
      {stage089[187]},
      {stage089[233]}
   );
   gpc1_1 gpc1_1_7015(
      {stage089[188]},
      {stage089[234]}
   );
   gpc1_1 gpc1_1_7016(
      {stage089[189]},
      {stage089[235]}
   );
   gpc1_1 gpc1_1_7017(
      {stage089[190]},
      {stage089[236]}
   );
   gpc1_1 gpc1_1_7018(
      {stage089[191]},
      {stage089[237]}
   );
   gpc1_1 gpc1_1_7019(
      {stage089[192]},
      {stage089[238]}
   );
   gpc1_1 gpc1_1_7020(
      {stage089[193]},
      {stage089[239]}
   );
   gpc1_1 gpc1_1_7021(
      {stage089[194]},
      {stage089[240]}
   );
   gpc1_1 gpc1_1_7022(
      {stage089[195]},
      {stage089[241]}
   );
   gpc1_1 gpc1_1_7023(
      {stage089[196]},
      {stage089[242]}
   );
   gpc1_1 gpc1_1_7024(
      {stage089[197]},
      {stage089[243]}
   );
   gpc606_5 gpc606_5_7025(
      {stage089[198], stage089[199], stage089[200], stage089[201], stage089[202], stage089[203]},
      {stage091[200], stage091[201], stage091[202], stage091[203], stage091[204], stage091[205]},
      {stage093[209], stage092[229], stage091[259], stage090[222], stage089[244]}
   );
   gpc606_5 gpc606_5_7026(
      {stage089[204], stage089[205], stage089[206], stage089[207], stage089[208], stage089[209]},
      {stage091[206], stage091[207], stage091[208], stage091[209], stage091[210], stage091[211]},
      {stage093[210], stage092[230], stage091[260], stage090[223], stage089[245]}
   );
   gpc606_5 gpc606_5_7027(
      {stage089[210], stage089[211], stage089[212], stage089[213], stage089[214], stage089[215]},
      {stage091[212], stage091[213], stage091[214], stage091[215], stage091[216], stage091[217]},
      {stage093[211], stage092[231], stage091[261], stage090[224], stage089[246]}
   );
   gpc1_1 gpc1_1_7028(
      {stage090[192]},
      {stage090[225]}
   );
   gpc1_1 gpc1_1_7029(
      {stage090[193]},
      {stage090[226]}
   );
   gpc606_5 gpc606_5_7030(
      {stage090[194], stage090[195], stage090[196], stage090[197], stage090[198], stage090[199]},
      {stage092[198], stage092[199], stage092[200], stage092[201], stage092[202], stage092[203]},
      {stage094[224], stage093[212], stage092[232], stage091[262], stage090[227]}
   );
   gpc606_5 gpc606_5_7031(
      {stage090[200], stage090[201], stage090[202], stage090[203], stage090[204], stage090[205]},
      {stage092[204], stage092[205], stage092[206], stage092[207], stage092[208], stage092[209]},
      {stage094[225], stage093[213], stage092[233], stage091[263], stage090[228]}
   );
   gpc606_5 gpc606_5_7032(
      {stage090[206], stage090[207], stage090[208], stage090[209], stage090[210], stage090[211]},
      {stage092[210], stage092[211], stage092[212], stage092[213], stage092[214], stage092[215]},
      {stage094[226], stage093[214], stage092[234], stage091[264], stage090[229]}
   );
   gpc615_5 gpc615_5_7033(
      {stage090[212], stage090[213], stage090[214], stage090[215], stage090[216]},
      {stage091[218]},
      {stage092[216], stage092[217], stage092[218], stage092[219], stage092[220], stage092[221]},
      {stage094[227], stage093[215], stage092[235], stage091[265], stage090[230]}
   );
   gpc1_1 gpc1_1_7034(
      {stage091[219]},
      {stage091[266]}
   );
   gpc1_1 gpc1_1_7035(
      {stage091[220]},
      {stage091[267]}
   );
   gpc1_1 gpc1_1_7036(
      {stage091[221]},
      {stage091[268]}
   );
   gpc1_1 gpc1_1_7037(
      {stage091[222]},
      {stage091[269]}
   );
   gpc1_1 gpc1_1_7038(
      {stage091[223]},
      {stage091[270]}
   );
   gpc1_1 gpc1_1_7039(
      {stage091[224]},
      {stage091[271]}
   );
   gpc1_1 gpc1_1_7040(
      {stage091[225]},
      {stage091[272]}
   );
   gpc1_1 gpc1_1_7041(
      {stage091[226]},
      {stage091[273]}
   );
   gpc1_1 gpc1_1_7042(
      {stage091[227]},
      {stage091[274]}
   );
   gpc1_1 gpc1_1_7043(
      {stage091[228]},
      {stage091[275]}
   );
   gpc1_1 gpc1_1_7044(
      {stage091[229]},
      {stage091[276]}
   );
   gpc1_1 gpc1_1_7045(
      {stage091[230]},
      {stage091[277]}
   );
   gpc1_1 gpc1_1_7046(
      {stage091[231]},
      {stage091[278]}
   );
   gpc1_1 gpc1_1_7047(
      {stage091[232]},
      {stage091[279]}
   );
   gpc1_1 gpc1_1_7048(
      {stage091[233]},
      {stage091[280]}
   );
   gpc1_1 gpc1_1_7049(
      {stage091[234]},
      {stage091[281]}
   );
   gpc1_1 gpc1_1_7050(
      {stage091[235]},
      {stage091[282]}
   );
   gpc1_1 gpc1_1_7051(
      {stage091[236]},
      {stage091[283]}
   );
   gpc1_1 gpc1_1_7052(
      {stage091[237]},
      {stage091[284]}
   );
   gpc1_1 gpc1_1_7053(
      {stage091[238]},
      {stage091[285]}
   );
   gpc1_1 gpc1_1_7054(
      {stage091[239]},
      {stage091[286]}
   );
   gpc1_1 gpc1_1_7055(
      {stage091[240]},
      {stage091[287]}
   );
   gpc1_1 gpc1_1_7056(
      {stage091[241]},
      {stage091[288]}
   );
   gpc1_1 gpc1_1_7057(
      {stage091[242]},
      {stage091[289]}
   );
   gpc1_1 gpc1_1_7058(
      {stage091[243]},
      {stage091[290]}
   );
   gpc1_1 gpc1_1_7059(
      {stage091[244]},
      {stage091[291]}
   );
   gpc1_1 gpc1_1_7060(
      {stage091[245]},
      {stage091[292]}
   );
   gpc1_1 gpc1_1_7061(
      {stage091[246]},
      {stage091[293]}
   );
   gpc1_1 gpc1_1_7062(
      {stage091[247]},
      {stage091[294]}
   );
   gpc1_1 gpc1_1_7063(
      {stage091[248]},
      {stage091[295]}
   );
   gpc1_1 gpc1_1_7064(
      {stage091[249]},
      {stage091[296]}
   );
   gpc1_1 gpc1_1_7065(
      {stage091[250]},
      {stage091[297]}
   );
   gpc1_1 gpc1_1_7066(
      {stage091[251]},
      {stage091[298]}
   );
   gpc1_1 gpc1_1_7067(
      {stage091[252]},
      {stage091[299]}
   );
   gpc1_1 gpc1_1_7068(
      {stage091[253]},
      {stage091[300]}
   );
   gpc1_1 gpc1_1_7069(
      {stage091[254]},
      {stage091[301]}
   );
   gpc1_1 gpc1_1_7070(
      {stage092[222]},
      {stage092[236]}
   );
   gpc1_1 gpc1_1_7071(
      {stage092[223]},
      {stage092[237]}
   );
   gpc1_1 gpc1_1_7072(
      {stage092[224]},
      {stage092[238]}
   );
   gpc1_1 gpc1_1_7073(
      {stage092[225]},
      {stage092[239]}
   );
   gpc1_1 gpc1_1_7074(
      {stage092[226]},
      {stage092[240]}
   );
   gpc1_1 gpc1_1_7075(
      {stage093[189]},
      {stage093[216]}
   );
   gpc1_1 gpc1_1_7076(
      {stage093[190]},
      {stage093[217]}
   );
   gpc606_5 gpc606_5_7077(
      {stage093[191], stage093[192], stage093[193], stage093[194], stage093[195], stage093[196]},
      {stage095[181], stage095[182], stage095[183], stage095[184], stage095[185], stage095[186]},
      {stage097[205], stage096[218], stage095[205], stage094[228], stage093[218]}
   );
   gpc606_5 gpc606_5_7078(
      {stage093[197], stage093[198], stage093[199], stage093[200], stage093[201], stage093[202]},
      {stage095[187], stage095[188], stage095[189], stage095[190], stage095[191], stage095[192]},
      {stage097[206], stage096[219], stage095[206], stage094[229], stage093[219]}
   );
   gpc606_5 gpc606_5_7079(
      {stage093[203], stage093[204], stage093[205], stage093[206], stage093[207], stage093[208]},
      {stage095[193], stage095[194], stage095[195], stage095[196], stage095[197], stage095[198]},
      {stage097[207], stage096[220], stage095[207], stage094[230], stage093[220]}
   );
   gpc606_5 gpc606_5_7080(
      {stage094[195], stage094[196], stage094[197], stage094[198], stage094[199], stage094[200]},
      {stage096[184], stage096[185], stage096[186], stage096[187], stage096[188], stage096[189]},
      {stage098[206], stage097[208], stage096[221], stage095[208], stage094[231]}
   );
   gpc606_5 gpc606_5_7081(
      {stage094[201], stage094[202], stage094[203], stage094[204], stage094[205], stage094[206]},
      {stage096[190], stage096[191], stage096[192], stage096[193], stage096[194], stage096[195]},
      {stage098[207], stage097[209], stage096[222], stage095[209], stage094[232]}
   );
   gpc606_5 gpc606_5_7082(
      {stage094[207], stage094[208], stage094[209], stage094[210], stage094[211], stage094[212]},
      {stage096[196], stage096[197], stage096[198], stage096[199], stage096[200], stage096[201]},
      {stage098[208], stage097[210], stage096[223], stage095[210], stage094[233]}
   );
   gpc606_5 gpc606_5_7083(
      {stage094[213], stage094[214], stage094[215], stage094[216], stage094[217], stage094[218]},
      {stage096[202], stage096[203], stage096[204], stage096[205], stage096[206], stage096[207]},
      {stage098[209], stage097[211], stage096[224], stage095[211], stage094[234]}
   );
   gpc606_5 gpc606_5_7084(
      {stage094[219], stage094[220], stage094[221], stage094[222], stage094[223], 1'h0},
      {stage096[208], stage096[209], stage096[210], stage096[211], stage096[212], stage096[213]},
      {stage098[210], stage097[212], stage096[225], stage095[212], stage094[235]}
   );
   gpc606_5 gpc606_5_7085(
      {stage095[199], stage095[200], stage095[201], stage095[202], stage095[203], stage095[204]},
      {stage097[175], stage097[176], stage097[177], stage097[178], stage097[179], stage097[180]},
      {stage099[258], stage098[211], stage097[213], stage096[226], stage095[213]}
   );
   gpc1_1 gpc1_1_7086(
      {stage096[214]},
      {stage096[227]}
   );
   gpc1_1 gpc1_1_7087(
      {stage096[215]},
      {stage096[228]}
   );
   gpc1_1 gpc1_1_7088(
      {stage096[216]},
      {stage096[229]}
   );
   gpc1_1 gpc1_1_7089(
      {stage096[217]},
      {stage096[230]}
   );
   gpc1_1 gpc1_1_7090(
      {stage097[181]},
      {stage097[214]}
   );
   gpc1_1 gpc1_1_7091(
      {stage097[182]},
      {stage097[215]}
   );
   gpc606_5 gpc606_5_7092(
      {stage097[183], stage097[184], stage097[185], stage097[186], stage097[187], stage097[188]},
      {stage099[204], stage099[205], stage099[206], stage099[207], stage099[208], stage099[209]},
      {stage101[229], stage100[202], stage099[259], stage098[212], stage097[216]}
   );
   gpc606_5 gpc606_5_7093(
      {stage097[189], stage097[190], stage097[191], stage097[192], stage097[193], stage097[194]},
      {stage099[210], stage099[211], stage099[212], stage099[213], stage099[214], stage099[215]},
      {stage101[230], stage100[203], stage099[260], stage098[213], stage097[217]}
   );
   gpc615_5 gpc615_5_7094(
      {stage097[195], stage097[196], stage097[197], stage097[198], stage097[199]},
      {stage098[184]},
      {stage099[216], stage099[217], stage099[218], stage099[219], stage099[220], stage099[221]},
      {stage101[231], stage100[204], stage099[261], stage098[214], stage097[218]}
   );
   gpc615_5 gpc615_5_7095(
      {stage097[200], stage097[201], stage097[202], stage097[203], stage097[204]},
      {stage098[185]},
      {stage099[222], stage099[223], stage099[224], stage099[225], stage099[226], stage099[227]},
      {stage101[232], stage100[205], stage099[262], stage098[215], stage097[219]}
   );
   gpc1_1 gpc1_1_7096(
      {stage098[186]},
      {stage098[216]}
   );
   gpc1_1 gpc1_1_7097(
      {stage098[187]},
      {stage098[217]}
   );
   gpc1_1 gpc1_1_7098(
      {stage098[188]},
      {stage098[218]}
   );
   gpc1_1 gpc1_1_7099(
      {stage098[189]},
      {stage098[219]}
   );
   gpc1_1 gpc1_1_7100(
      {stage098[190]},
      {stage098[220]}
   );
   gpc1_1 gpc1_1_7101(
      {stage098[191]},
      {stage098[221]}
   );
   gpc1_1 gpc1_1_7102(
      {stage098[192]},
      {stage098[222]}
   );
   gpc1_1 gpc1_1_7103(
      {stage098[193]},
      {stage098[223]}
   );
   gpc606_5 gpc606_5_7104(
      {stage098[194], stage098[195], stage098[196], stage098[197], stage098[198], stage098[199]},
      {stage100[178], stage100[179], stage100[180], stage100[181], stage100[182], stage100[183]},
      {stage102[221], stage101[233], stage100[206], stage099[263], stage098[224]}
   );
   gpc606_5 gpc606_5_7105(
      {stage098[200], stage098[201], stage098[202], stage098[203], stage098[204], stage098[205]},
      {stage100[184], stage100[185], stage100[186], stage100[187], stage100[188], stage100[189]},
      {stage102[222], stage101[234], stage100[207], stage099[264], stage098[225]}
   );
   gpc1_1 gpc1_1_7106(
      {stage099[228]},
      {stage099[265]}
   );
   gpc1_1 gpc1_1_7107(
      {stage099[229]},
      {stage099[266]}
   );
   gpc1_1 gpc1_1_7108(
      {stage099[230]},
      {stage099[267]}
   );
   gpc1_1 gpc1_1_7109(
      {stage099[231]},
      {stage099[268]}
   );
   gpc1_1 gpc1_1_7110(
      {stage099[232]},
      {stage099[269]}
   );
   gpc1_1 gpc1_1_7111(
      {stage099[233]},
      {stage099[270]}
   );
   gpc1_1 gpc1_1_7112(
      {stage099[234]},
      {stage099[271]}
   );
   gpc1_1 gpc1_1_7113(
      {stage099[235]},
      {stage099[272]}
   );
   gpc1_1 gpc1_1_7114(
      {stage099[236]},
      {stage099[273]}
   );
   gpc1_1 gpc1_1_7115(
      {stage099[237]},
      {stage099[274]}
   );
   gpc1_1 gpc1_1_7116(
      {stage099[238]},
      {stage099[275]}
   );
   gpc1_1 gpc1_1_7117(
      {stage099[239]},
      {stage099[276]}
   );
   gpc606_5 gpc606_5_7118(
      {stage099[240], stage099[241], stage099[242], stage099[243], stage099[244], stage099[245]},
      {stage101[192], stage101[193], stage101[194], stage101[195], stage101[196], stage101[197]},
      {stage103[225], stage102[223], stage101[235], stage100[208], stage099[277]}
   );
   gpc606_5 gpc606_5_7119(
      {stage099[246], stage099[247], stage099[248], stage099[249], stage099[250], stage099[251]},
      {stage101[198], stage101[199], stage101[200], stage101[201], stage101[202], stage101[203]},
      {stage103[226], stage102[224], stage101[236], stage100[209], stage099[278]}
   );
   gpc606_5 gpc606_5_7120(
      {stage099[252], stage099[253], stage099[254], stage099[255], stage099[256], stage099[257]},
      {stage101[204], stage101[205], stage101[206], stage101[207], stage101[208], stage101[209]},
      {stage103[227], stage102[225], stage101[237], stage100[210], stage099[279]}
   );
   gpc1_1 gpc1_1_7121(
      {stage100[190]},
      {stage100[211]}
   );
   gpc1_1 gpc1_1_7122(
      {stage100[191]},
      {stage100[212]}
   );
   gpc1_1 gpc1_1_7123(
      {stage100[192]},
      {stage100[213]}
   );
   gpc1_1 gpc1_1_7124(
      {stage100[193]},
      {stage100[214]}
   );
   gpc1_1 gpc1_1_7125(
      {stage100[194]},
      {stage100[215]}
   );
   gpc1_1 gpc1_1_7126(
      {stage100[195]},
      {stage100[216]}
   );
   gpc1406_5 gpc1406_5_7127(
      {stage100[196], stage100[197], stage100[198], stage100[199], stage100[200], stage100[201]},
      {stage102[200], stage102[201], stage102[202], stage102[203]},
      {stage103[192]},
      {stage104[245], stage103[228], stage102[226], stage101[238], stage100[217]}
   );
   gpc1_1 gpc1_1_7128(
      {stage101[210]},
      {stage101[239]}
   );
   gpc1_1 gpc1_1_7129(
      {stage101[211]},
      {stage101[240]}
   );
   gpc1_1 gpc1_1_7130(
      {stage101[212]},
      {stage101[241]}
   );
   gpc1_1 gpc1_1_7131(
      {stage101[213]},
      {stage101[242]}
   );
   gpc1_1 gpc1_1_7132(
      {stage101[214]},
      {stage101[243]}
   );
   gpc1_1 gpc1_1_7133(
      {stage101[215]},
      {stage101[244]}
   );
   gpc1_1 gpc1_1_7134(
      {stage101[216]},
      {stage101[245]}
   );
   gpc1_1 gpc1_1_7135(
      {stage101[217]},
      {stage101[246]}
   );
   gpc1_1 gpc1_1_7136(
      {stage101[218]},
      {stage101[247]}
   );
   gpc1_1 gpc1_1_7137(
      {stage101[219]},
      {stage101[248]}
   );
   gpc1_1 gpc1_1_7138(
      {stage101[220]},
      {stage101[249]}
   );
   gpc1_1 gpc1_1_7139(
      {stage101[221]},
      {stage101[250]}
   );
   gpc1_1 gpc1_1_7140(
      {stage101[222]},
      {stage101[251]}
   );
   gpc606_5 gpc606_5_7141(
      {stage101[223], stage101[224], stage101[225], stage101[226], stage101[227], stage101[228]},
      {stage103[193], stage103[194], stage103[195], stage103[196], stage103[197], stage103[198]},
      {stage105[206], stage104[246], stage103[229], stage102[227], stage101[252]}
   );
   gpc1_1 gpc1_1_7142(
      {stage102[204]},
      {stage102[228]}
   );
   gpc1_1 gpc1_1_7143(
      {stage102[205]},
      {stage102[229]}
   );
   gpc1_1 gpc1_1_7144(
      {stage102[206]},
      {stage102[230]}
   );
   gpc623_5 gpc623_5_7145(
      {stage102[207], stage102[208], stage102[209]},
      {stage103[199], stage103[200]},
      {stage104[211], stage104[212], stage104[213], stage104[214], stage104[215], stage104[216]},
      {stage106[229], stage105[207], stage104[247], stage103[230], stage102[231]}
   );
   gpc615_5 gpc615_5_7146(
      {stage102[210], stage102[211], stage102[212], stage102[213], stage102[214]},
      {stage103[201]},
      {stage104[217], stage104[218], stage104[219], stage104[220], stage104[221], stage104[222]},
      {stage106[230], stage105[208], stage104[248], stage103[231], stage102[232]}
   );
   gpc1343_5 gpc1343_5_7147(
      {stage102[215], stage102[216], stage102[217]},
      {stage103[202], stage103[203], stage103[204], stage103[205]},
      {stage104[223], stage104[224], stage104[225]},
      {stage105[183]},
      {stage106[231], stage105[209], stage104[249], stage103[232], stage102[233]}
   );
   gpc1343_5 gpc1343_5_7148(
      {stage102[218], stage102[219], stage102[220]},
      {stage103[206], stage103[207], stage103[208], stage103[209]},
      {stage104[226], stage104[227], stage104[228]},
      {stage105[184]},
      {stage106[232], stage105[210], stage104[250], stage103[233], stage102[234]}
   );
   gpc615_5 gpc615_5_7149(
      {stage103[210], stage103[211], stage103[212], stage103[213], stage103[214]},
      {stage104[229]},
      {stage105[185], stage105[186], stage105[187], stage105[188], stage105[189], stage105[190]},
      {stage107[228], stage106[233], stage105[211], stage104[251], stage103[234]}
   );
   gpc615_5 gpc615_5_7150(
      {stage103[215], stage103[216], stage103[217], stage103[218], stage103[219]},
      {stage104[230]},
      {stage105[191], stage105[192], stage105[193], stage105[194], stage105[195], stage105[196]},
      {stage107[229], stage106[234], stage105[212], stage104[252], stage103[235]}
   );
   gpc615_5 gpc615_5_7151(
      {stage103[220], stage103[221], stage103[222], stage103[223], stage103[224]},
      {stage104[231]},
      {stage105[197], stage105[198], stage105[199], stage105[200], stage105[201], stage105[202]},
      {stage107[230], stage106[235], stage105[213], stage104[253], stage103[236]}
   );
   gpc1_1 gpc1_1_7152(
      {stage104[232]},
      {stage104[254]}
   );
   gpc606_5 gpc606_5_7153(
      {stage104[233], stage104[234], stage104[235], stage104[236], stage104[237], stage104[238]},
      {stage106[197], stage106[198], stage106[199], stage106[200], stage106[201], stage106[202]},
      {stage108[225], stage107[231], stage106[236], stage105[214], stage104[255]}
   );
   gpc606_5 gpc606_5_7154(
      {stage104[239], stage104[240], stage104[241], stage104[242], stage104[243], stage104[244]},
      {stage106[203], stage106[204], stage106[205], stage106[206], stage106[207], stage106[208]},
      {stage108[226], stage107[232], stage106[237], stage105[215], stage104[256]}
   );
   gpc615_5 gpc615_5_7155(
      {stage105[203], stage105[204], stage105[205], 1'h0, 1'h0},
      {stage106[209]},
      {stage107[187], stage107[188], stage107[189], stage107[190], stage107[191], stage107[192]},
      {stage109[209], stage108[227], stage107[233], stage106[238], stage105[216]}
   );
   gpc1_1 gpc1_1_7156(
      {stage106[210]},
      {stage106[239]}
   );
   gpc1_1 gpc1_1_7157(
      {stage106[211]},
      {stage106[240]}
   );
   gpc1_1 gpc1_1_7158(
      {stage106[212]},
      {stage106[241]}
   );
   gpc1_1 gpc1_1_7159(
      {stage106[213]},
      {stage106[242]}
   );
   gpc1_1 gpc1_1_7160(
      {stage106[214]},
      {stage106[243]}
   );
   gpc1_1 gpc1_1_7161(
      {stage106[215]},
      {stage106[244]}
   );
   gpc1_1 gpc1_1_7162(
      {stage106[216]},
      {stage106[245]}
   );
   gpc606_5 gpc606_5_7163(
      {stage106[217], stage106[218], stage106[219], stage106[220], stage106[221], stage106[222]},
      {stage108[180], stage108[181], stage108[182], stage108[183], stage108[184], stage108[185]},
      {stage110[236], stage109[210], stage108[228], stage107[234], stage106[246]}
   );
   gpc606_5 gpc606_5_7164(
      {stage106[223], stage106[224], stage106[225], stage106[226], stage106[227], stage106[228]},
      {stage108[186], stage108[187], stage108[188], stage108[189], stage108[190], stage108[191]},
      {stage110[237], stage109[211], stage108[229], stage107[235], stage106[247]}
   );
   gpc1_1 gpc1_1_7165(
      {stage107[193]},
      {stage107[236]}
   );
   gpc1_1 gpc1_1_7166(
      {stage107[194]},
      {stage107[237]}
   );
   gpc1_1 gpc1_1_7167(
      {stage107[195]},
      {stage107[238]}
   );
   gpc1_1 gpc1_1_7168(
      {stage107[196]},
      {stage107[239]}
   );
   gpc1_1 gpc1_1_7169(
      {stage107[197]},
      {stage107[240]}
   );
   gpc1_1 gpc1_1_7170(
      {stage107[198]},
      {stage107[241]}
   );
   gpc1_1 gpc1_1_7171(
      {stage107[199]},
      {stage107[242]}
   );
   gpc1_1 gpc1_1_7172(
      {stage107[200]},
      {stage107[243]}
   );
   gpc7_3 gpc7_3_7173(
      {stage107[201], stage107[202], stage107[203], stage107[204], stage107[205], stage107[206], stage107[207]},
      {stage109[212], stage108[230], stage107[244]}
   );
   gpc7_3 gpc7_3_7174(
      {stage107[208], stage107[209], stage107[210], stage107[211], stage107[212], stage107[213], stage107[214]},
      {stage109[213], stage108[231], stage107[245]}
   );
   gpc7_3 gpc7_3_7175(
      {stage107[215], stage107[216], stage107[217], stage107[218], stage107[219], stage107[220], stage107[221]},
      {stage109[214], stage108[232], stage107[246]}
   );
   gpc606_5 gpc606_5_7176(
      {stage107[222], stage107[223], stage107[224], stage107[225], stage107[226], stage107[227]},
      {stage109[183], stage109[184], stage109[185], stage109[186], stage109[187], stage109[188]},
      {stage111[242], stage110[238], stage109[215], stage108[233], stage107[247]}
   );
   gpc1_1 gpc1_1_7177(
      {stage108[192]},
      {stage108[234]}
   );
   gpc1_1 gpc1_1_7178(
      {stage108[193]},
      {stage108[235]}
   );
   gpc1_1 gpc1_1_7179(
      {stage108[194]},
      {stage108[236]}
   );
   gpc1_1 gpc1_1_7180(
      {stage108[195]},
      {stage108[237]}
   );
   gpc1_1 gpc1_1_7181(
      {stage108[196]},
      {stage108[238]}
   );
   gpc1_1 gpc1_1_7182(
      {stage108[197]},
      {stage108[239]}
   );
   gpc1_1 gpc1_1_7183(
      {stage108[198]},
      {stage108[240]}
   );
   gpc1_1 gpc1_1_7184(
      {stage108[199]},
      {stage108[241]}
   );
   gpc1_1 gpc1_1_7185(
      {stage108[200]},
      {stage108[242]}
   );
   gpc606_5 gpc606_5_7186(
      {stage108[201], stage108[202], stage108[203], stage108[204], stage108[205], stage108[206]},
      {stage110[199], stage110[200], stage110[201], stage110[202], stage110[203], stage110[204]},
      {stage112[215], stage111[243], stage110[239], stage109[216], stage108[243]}
   );
   gpc606_5 gpc606_5_7187(
      {stage108[207], stage108[208], stage108[209], stage108[210], stage108[211], stage108[212]},
      {stage110[205], stage110[206], stage110[207], stage110[208], stage110[209], stage110[210]},
      {stage112[216], stage111[244], stage110[240], stage109[217], stage108[244]}
   );
   gpc606_5 gpc606_5_7188(
      {stage108[213], stage108[214], stage108[215], stage108[216], stage108[217], stage108[218]},
      {stage110[211], stage110[212], stage110[213], stage110[214], stage110[215], stage110[216]},
      {stage112[217], stage111[245], stage110[241], stage109[218], stage108[245]}
   );
   gpc606_5 gpc606_5_7189(
      {stage108[219], stage108[220], stage108[221], stage108[222], stage108[223], stage108[224]},
      {stage110[217], stage110[218], stage110[219], stage110[220], stage110[221], stage110[222]},
      {stage112[218], stage111[246], stage110[242], stage109[219], stage108[246]}
   );
   gpc615_5 gpc615_5_7190(
      {stage109[189], stage109[190], stage109[191], stage109[192], stage109[193]},
      {stage110[223]},
      {stage111[215], stage111[216], stage111[217], stage111[218], stage111[219], stage111[220]},
      {stage113[213], stage112[219], stage111[247], stage110[243], stage109[220]}
   );
   gpc615_5 gpc615_5_7191(
      {stage109[194], stage109[195], stage109[196], stage109[197], stage109[198]},
      {stage110[224]},
      {stage111[221], stage111[222], stage111[223], stage111[224], stage111[225], stage111[226]},
      {stage113[214], stage112[220], stage111[248], stage110[244], stage109[221]}
   );
   gpc615_5 gpc615_5_7192(
      {stage109[199], stage109[200], stage109[201], stage109[202], stage109[203]},
      {stage110[225]},
      {stage111[227], stage111[228], stage111[229], stage111[230], stage111[231], stage111[232]},
      {stage113[215], stage112[221], stage111[249], stage110[245], stage109[222]}
   );
   gpc615_5 gpc615_5_7193(
      {stage109[204], stage109[205], stage109[206], stage109[207], stage109[208]},
      {stage110[226]},
      {stage111[233], stage111[234], stage111[235], stage111[236], stage111[237], stage111[238]},
      {stage113[216], stage112[222], stage111[250], stage110[246], stage109[223]}
   );
   gpc1_1 gpc1_1_7194(
      {stage110[227]},
      {stage110[247]}
   );
   gpc1_1 gpc1_1_7195(
      {stage110[228]},
      {stage110[248]}
   );
   gpc1_1 gpc1_1_7196(
      {stage110[229]},
      {stage110[249]}
   );
   gpc1_1 gpc1_1_7197(
      {stage110[230]},
      {stage110[250]}
   );
   gpc1_1 gpc1_1_7198(
      {stage110[231]},
      {stage110[251]}
   );
   gpc1_1 gpc1_1_7199(
      {stage110[232]},
      {stage110[252]}
   );
   gpc1_1 gpc1_1_7200(
      {stage110[233]},
      {stage110[253]}
   );
   gpc1_1 gpc1_1_7201(
      {stage110[234]},
      {stage110[254]}
   );
   gpc1_1 gpc1_1_7202(
      {stage110[235]},
      {stage110[255]}
   );
   gpc1_1 gpc1_1_7203(
      {stage111[239]},
      {stage111[251]}
   );
   gpc1_1 gpc1_1_7204(
      {stage111[240]},
      {stage111[252]}
   );
   gpc1_1 gpc1_1_7205(
      {stage111[241]},
      {stage111[253]}
   );
   gpc606_5 gpc606_5_7206(
      {stage112[192], stage112[193], stage112[194], stage112[195], stage112[196], stage112[197]},
      {stage114[183], stage114[184], stage114[185], stage114[186], stage114[187], stage114[188]},
      {stage116[214], stage115[237], stage114[216], stage113[217], stage112[223]}
   );
   gpc606_5 gpc606_5_7207(
      {stage112[198], stage112[199], stage112[200], stage112[201], stage112[202], stage112[203]},
      {stage114[189], stage114[190], stage114[191], stage114[192], stage114[193], stage114[194]},
      {stage116[215], stage115[238], stage114[217], stage113[218], stage112[224]}
   );
   gpc606_5 gpc606_5_7208(
      {stage112[204], stage112[205], stage112[206], stage112[207], stage112[208], stage112[209]},
      {stage114[195], stage114[196], stage114[197], stage114[198], stage114[199], stage114[200]},
      {stage116[216], stage115[239], stage114[218], stage113[219], stage112[225]}
   );
   gpc606_5 gpc606_5_7209(
      {stage112[210], stage112[211], stage112[212], stage112[213], stage112[214], 1'h0},
      {stage114[201], stage114[202], stage114[203], stage114[204], stage114[205], stage114[206]},
      {stage116[217], stage115[240], stage114[219], stage113[220], stage112[226]}
   );
   gpc606_5 gpc606_5_7210(
      {stage113[183], stage113[184], stage113[185], stage113[186], stage113[187], stage113[188]},
      {stage115[196], stage115[197], stage115[198], stage115[199], stage115[200], stage115[201]},
      {stage117[223], stage116[218], stage115[241], stage114[220], stage113[221]}
   );
   gpc606_5 gpc606_5_7211(
      {stage113[189], stage113[190], stage113[191], stage113[192], stage113[193], stage113[194]},
      {stage115[202], stage115[203], stage115[204], stage115[205], stage115[206], stage115[207]},
      {stage117[224], stage116[219], stage115[242], stage114[221], stage113[222]}
   );
   gpc606_5 gpc606_5_7212(
      {stage113[195], stage113[196], stage113[197], stage113[198], stage113[199], stage113[200]},
      {stage115[208], stage115[209], stage115[210], stage115[211], stage115[212], stage115[213]},
      {stage117[225], stage116[220], stage115[243], stage114[222], stage113[223]}
   );
   gpc606_5 gpc606_5_7213(
      {stage113[201], stage113[202], stage113[203], stage113[204], stage113[205], stage113[206]},
      {stage115[214], stage115[215], stage115[216], stage115[217], stage115[218], stage115[219]},
      {stage117[226], stage116[221], stage115[244], stage114[223], stage113[224]}
   );
   gpc606_5 gpc606_5_7214(
      {stage113[207], stage113[208], stage113[209], stage113[210], stage113[211], stage113[212]},
      {stage115[220], stage115[221], stage115[222], stage115[223], stage115[224], stage115[225]},
      {stage117[227], stage116[222], stage115[245], stage114[224], stage113[225]}
   );
   gpc1_1 gpc1_1_7215(
      {stage114[207]},
      {stage114[225]}
   );
   gpc1_1 gpc1_1_7216(
      {stage114[208]},
      {stage114[226]}
   );
   gpc1_1 gpc1_1_7217(
      {stage114[209]},
      {stage114[227]}
   );
   gpc1_1 gpc1_1_7218(
      {stage114[210]},
      {stage114[228]}
   );
   gpc1_1 gpc1_1_7219(
      {stage114[211]},
      {stage114[229]}
   );
   gpc1_1 gpc1_1_7220(
      {stage114[212]},
      {stage114[230]}
   );
   gpc1_1 gpc1_1_7221(
      {stage114[213]},
      {stage114[231]}
   );
   gpc1_1 gpc1_1_7222(
      {stage114[214]},
      {stage114[232]}
   );
   gpc1_1 gpc1_1_7223(
      {stage114[215]},
      {stage114[233]}
   );
   gpc1_1 gpc1_1_7224(
      {stage115[226]},
      {stage115[246]}
   );
   gpc1_1 gpc1_1_7225(
      {stage115[227]},
      {stage115[247]}
   );
   gpc1_1 gpc1_1_7226(
      {stage115[228]},
      {stage115[248]}
   );
   gpc1_1 gpc1_1_7227(
      {stage115[229]},
      {stage115[249]}
   );
   gpc1_1 gpc1_1_7228(
      {stage115[230]},
      {stage115[250]}
   );
   gpc606_5 gpc606_5_7229(
      {stage115[231], stage115[232], stage115[233], stage115[234], stage115[235], stage115[236]},
      {stage117[196], stage117[197], stage117[198], stage117[199], stage117[200], stage117[201]},
      {stage119[210], stage118[224], stage117[228], stage116[223], stage115[251]}
   );
   gpc1_1 gpc1_1_7230(
      {stage116[187]},
      {stage116[224]}
   );
   gpc1_1 gpc1_1_7231(
      {stage116[188]},
      {stage116[225]}
   );
   gpc1_1 gpc1_1_7232(
      {stage116[189]},
      {stage116[226]}
   );
   gpc606_5 gpc606_5_7233(
      {stage116[190], stage116[191], stage116[192], stage116[193], stage116[194], stage116[195]},
      {stage118[183], stage118[184], stage118[185], stage118[186], stage118[187], stage118[188]},
      {stage120[220], stage119[211], stage118[225], stage117[229], stage116[227]}
   );
   gpc606_5 gpc606_5_7234(
      {stage116[196], stage116[197], stage116[198], stage116[199], stage116[200], stage116[201]},
      {stage118[189], stage118[190], stage118[191], stage118[192], stage118[193], stage118[194]},
      {stage120[221], stage119[212], stage118[226], stage117[230], stage116[228]}
   );
   gpc606_5 gpc606_5_7235(
      {stage116[202], stage116[203], stage116[204], stage116[205], stage116[206], stage116[207]},
      {stage118[195], stage118[196], stage118[197], stage118[198], stage118[199], stage118[200]},
      {stage120[222], stage119[213], stage118[227], stage117[231], stage116[229]}
   );
   gpc606_5 gpc606_5_7236(
      {stage116[208], stage116[209], stage116[210], stage116[211], stage116[212], stage116[213]},
      {stage118[201], stage118[202], stage118[203], stage118[204], stage118[205], stage118[206]},
      {stage120[223], stage119[214], stage118[228], stage117[232], stage116[230]}
   );
   gpc1_1 gpc1_1_7237(
      {stage117[202]},
      {stage117[233]}
   );
   gpc1_1 gpc1_1_7238(
      {stage117[203]},
      {stage117[234]}
   );
   gpc1_1 gpc1_1_7239(
      {stage117[204]},
      {stage117[235]}
   );
   gpc1_1 gpc1_1_7240(
      {stage117[205]},
      {stage117[236]}
   );
   gpc1_1 gpc1_1_7241(
      {stage117[206]},
      {stage117[237]}
   );
   gpc1_1 gpc1_1_7242(
      {stage117[207]},
      {stage117[238]}
   );
   gpc1_1 gpc1_1_7243(
      {stage117[208]},
      {stage117[239]}
   );
   gpc1_1 gpc1_1_7244(
      {stage117[209]},
      {stage117[240]}
   );
   gpc1_1 gpc1_1_7245(
      {stage117[210]},
      {stage117[241]}
   );
   gpc606_5 gpc606_5_7246(
      {stage117[211], stage117[212], stage117[213], stage117[214], stage117[215], stage117[216]},
      {stage119[184], stage119[185], stage119[186], stage119[187], stage119[188], stage119[189]},
      {stage121[205], stage120[224], stage119[215], stage118[229], stage117[242]}
   );
   gpc606_5 gpc606_5_7247(
      {stage117[217], stage117[218], stage117[219], stage117[220], stage117[221], stage117[222]},
      {stage119[190], stage119[191], stage119[192], stage119[193], stage119[194], stage119[195]},
      {stage121[206], stage120[225], stage119[216], stage118[230], stage117[243]}
   );
   gpc1_1 gpc1_1_7248(
      {stage118[207]},
      {stage118[231]}
   );
   gpc1_1 gpc1_1_7249(
      {stage118[208]},
      {stage118[232]}
   );
   gpc1_1 gpc1_1_7250(
      {stage118[209]},
      {stage118[233]}
   );
   gpc1_1 gpc1_1_7251(
      {stage118[210]},
      {stage118[234]}
   );
   gpc1_1 gpc1_1_7252(
      {stage118[211]},
      {stage118[235]}
   );
   gpc1_1 gpc1_1_7253(
      {stage118[212]},
      {stage118[236]}
   );
   gpc1_1 gpc1_1_7254(
      {stage118[213]},
      {stage118[237]}
   );
   gpc1_1 gpc1_1_7255(
      {stage118[214]},
      {stage118[238]}
   );
   gpc1_1 gpc1_1_7256(
      {stage118[215]},
      {stage118[239]}
   );
   gpc1_1 gpc1_1_7257(
      {stage118[216]},
      {stage118[240]}
   );
   gpc1_1 gpc1_1_7258(
      {stage118[217]},
      {stage118[241]}
   );
   gpc1_1 gpc1_1_7259(
      {stage118[218]},
      {stage118[242]}
   );
   gpc1_1 gpc1_1_7260(
      {stage118[219]},
      {stage118[243]}
   );
   gpc1_1 gpc1_1_7261(
      {stage118[220]},
      {stage118[244]}
   );
   gpc1_1 gpc1_1_7262(
      {stage118[221]},
      {stage118[245]}
   );
   gpc1_1 gpc1_1_7263(
      {stage118[222]},
      {stage118[246]}
   );
   gpc1_1 gpc1_1_7264(
      {stage118[223]},
      {stage118[247]}
   );
   gpc606_5 gpc606_5_7265(
      {stage119[196], stage119[197], stage119[198], stage119[199], stage119[200], stage119[201]},
      {stage121[176], stage121[177], stage121[178], stage121[179], stage121[180], stage121[181]},
      {stage123[282], stage122[222], stage121[207], stage120[226], stage119[217]}
   );
   gpc606_5 gpc606_5_7266(
      {stage119[202], stage119[203], stage119[204], stage119[205], stage119[206], stage119[207]},
      {stage121[182], stage121[183], stage121[184], stage121[185], stage121[186], stage121[187]},
      {stage123[283], stage122[223], stage121[208], stage120[227], stage119[218]}
   );
   gpc606_5 gpc606_5_7267(
      {stage119[208], stage119[209], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage121[188], stage121[189], stage121[190], stage121[191], stage121[192], stage121[193]},
      {stage123[284], stage122[224], stage121[209], stage120[228], stage119[219]}
   );
   gpc1_1 gpc1_1_7268(
      {stage120[185]},
      {stage120[229]}
   );
   gpc1_1 gpc1_1_7269(
      {stage120[186]},
      {stage120[230]}
   );
   gpc1_1 gpc1_1_7270(
      {stage120[187]},
      {stage120[231]}
   );
   gpc1_1 gpc1_1_7271(
      {stage120[188]},
      {stage120[232]}
   );
   gpc1_1 gpc1_1_7272(
      {stage120[189]},
      {stage120[233]}
   );
   gpc1_1 gpc1_1_7273(
      {stage120[190]},
      {stage120[234]}
   );
   gpc1_1 gpc1_1_7274(
      {stage120[191]},
      {stage120[235]}
   );
   gpc1_1 gpc1_1_7275(
      {stage120[192]},
      {stage120[236]}
   );
   gpc1_1 gpc1_1_7276(
      {stage120[193]},
      {stage120[237]}
   );
   gpc1_1 gpc1_1_7277(
      {stage120[194]},
      {stage120[238]}
   );
   gpc1_1 gpc1_1_7278(
      {stage120[195]},
      {stage120[239]}
   );
   gpc1_1 gpc1_1_7279(
      {stage120[196]},
      {stage120[240]}
   );
   gpc606_5 gpc606_5_7280(
      {stage120[197], stage120[198], stage120[199], stage120[200], stage120[201], stage120[202]},
      {stage122[187], stage122[188], stage122[189], stage122[190], stage122[191], stage122[192]},
      {stage124[212], stage123[285], stage122[225], stage121[210], stage120[241]}
   );
   gpc606_5 gpc606_5_7281(
      {stage120[203], stage120[204], stage120[205], stage120[206], stage120[207], stage120[208]},
      {stage122[193], stage122[194], stage122[195], stage122[196], stage122[197], stage122[198]},
      {stage124[213], stage123[286], stage122[226], stage121[211], stage120[242]}
   );
   gpc606_5 gpc606_5_7282(
      {stage120[209], stage120[210], stage120[211], stage120[212], stage120[213], stage120[214]},
      {stage122[199], stage122[200], stage122[201], stage122[202], stage122[203], stage122[204]},
      {stage124[214], stage123[287], stage122[227], stage121[212], stage120[243]}
   );
   gpc615_5 gpc615_5_7283(
      {stage120[215], stage120[216], stage120[217], stage120[218], stage120[219]},
      {stage121[194]},
      {stage122[205], stage122[206], stage122[207], stage122[208], stage122[209], stage122[210]},
      {stage124[215], stage123[288], stage122[228], stage121[213], stage120[244]}
   );
   gpc1_1 gpc1_1_7284(
      {stage121[195]},
      {stage121[214]}
   );
   gpc623_5 gpc623_5_7285(
      {stage121[196], stage121[197], stage121[198]},
      {stage122[211], stage122[212]},
      {stage123[256], stage123[257], stage123[258], stage123[259], stage123[260], stage123[261]},
      {stage125[241], stage124[216], stage123[289], stage122[229], stage121[215]}
   );
   gpc606_5 gpc606_5_7286(
      {stage121[199], stage121[200], stage121[201], stage121[202], stage121[203], stage121[204]},
      {stage123[262], stage123[263], stage123[264], stage123[265], stage123[266], stage123[267]},
      {stage125[242], stage124[217], stage123[290], stage122[230], stage121[216]}
   );
   gpc1_1 gpc1_1_7287(
      {stage122[213]},
      {stage122[231]}
   );
   gpc1_1 gpc1_1_7288(
      {stage122[214]},
      {stage122[232]}
   );
   gpc1_1 gpc1_1_7289(
      {stage122[215]},
      {stage122[233]}
   );
   gpc606_5 gpc606_5_7290(
      {stage122[216], stage122[217], stage122[218], stage122[219], stage122[220], stage122[221]},
      {stage124[178], stage124[179], stage124[180], stage124[181], stage124[182], stage124[183]},
      {stage126[242], stage125[243], stage124[218], stage123[291], stage122[234]}
   );
   gpc1_1 gpc1_1_7291(
      {stage123[268]},
      {stage123[292]}
   );
   gpc1_1 gpc1_1_7292(
      {stage123[269]},
      {stage123[293]}
   );
   gpc1_1 gpc1_1_7293(
      {stage123[270]},
      {stage123[294]}
   );
   gpc1_1 gpc1_1_7294(
      {stage123[271]},
      {stage123[295]}
   );
   gpc1_1 gpc1_1_7295(
      {stage123[272]},
      {stage123[296]}
   );
   gpc1_1 gpc1_1_7296(
      {stage123[273]},
      {stage123[297]}
   );
   gpc1_1 gpc1_1_7297(
      {stage123[274]},
      {stage123[298]}
   );
   gpc1_1 gpc1_1_7298(
      {stage123[275]},
      {stage123[299]}
   );
   gpc1_1 gpc1_1_7299(
      {stage123[276]},
      {stage123[300]}
   );
   gpc1_1 gpc1_1_7300(
      {stage123[277]},
      {stage123[301]}
   );
   gpc1_1 gpc1_1_7301(
      {stage123[278]},
      {stage123[302]}
   );
   gpc1_1 gpc1_1_7302(
      {stage123[279]},
      {stage123[303]}
   );
   gpc1_1 gpc1_1_7303(
      {stage123[280]},
      {stage123[304]}
   );
   gpc1_1 gpc1_1_7304(
      {stage123[281]},
      {stage123[305]}
   );
   gpc606_5 gpc606_5_7305(
      {stage124[184], stage124[185], stage124[186], stage124[187], stage124[188], stage124[189]},
      {stage126[189], stage126[190], stage126[191], stage126[192], stage126[193], stage126[194]},
      {stage128[47], stage127[254], stage126[243], stage125[244], stage124[219]}
   );
   gpc606_5 gpc606_5_7306(
      {stage124[190], stage124[191], stage124[192], stage124[193], stage124[194], stage124[195]},
      {stage126[195], stage126[196], stage126[197], stage126[198], stage126[199], stage126[200]},
      {stage128[48], stage127[255], stage126[244], stage125[245], stage124[220]}
   );
   gpc606_5 gpc606_5_7307(
      {stage124[196], stage124[197], stage124[198], stage124[199], stage124[200], stage124[201]},
      {stage126[201], stage126[202], stage126[203], stage126[204], stage126[205], stage126[206]},
      {stage128[49], stage127[256], stage126[245], stage125[246], stage124[221]}
   );
   gpc615_5 gpc615_5_7308(
      {stage124[202], stage124[203], stage124[204], stage124[205], stage124[206]},
      {stage125[205]},
      {stage126[207], stage126[208], stage126[209], stage126[210], stage126[211], stage126[212]},
      {stage128[50], stage127[257], stage126[246], stage125[247], stage124[222]}
   );
   gpc615_5 gpc615_5_7309(
      {stage124[207], stage124[208], stage124[209], stage124[210], stage124[211]},
      {stage125[206]},
      {stage126[213], stage126[214], stage126[215], stage126[216], stage126[217], stage126[218]},
      {stage128[51], stage127[258], stage126[247], stage125[248], stage124[223]}
   );
   gpc1_1 gpc1_1_7310(
      {stage125[207]},
      {stage125[249]}
   );
   gpc1_1 gpc1_1_7311(
      {stage125[208]},
      {stage125[250]}
   );
   gpc1_1 gpc1_1_7312(
      {stage125[209]},
      {stage125[251]}
   );
   gpc1_1 gpc1_1_7313(
      {stage125[210]},
      {stage125[252]}
   );
   gpc1_1 gpc1_1_7314(
      {stage125[211]},
      {stage125[253]}
   );
   gpc1_1 gpc1_1_7315(
      {stage125[212]},
      {stage125[254]}
   );
   gpc1_1 gpc1_1_7316(
      {stage125[213]},
      {stage125[255]}
   );
   gpc1_1 gpc1_1_7317(
      {stage125[214]},
      {stage125[256]}
   );
   gpc1_1 gpc1_1_7318(
      {stage125[215]},
      {stage125[257]}
   );
   gpc1_1 gpc1_1_7319(
      {stage125[216]},
      {stage125[258]}
   );
   gpc606_5 gpc606_5_7320(
      {stage125[217], stage125[218], stage125[219], stage125[220], stage125[221], stage125[222]},
      {stage127[212], stage127[213], stage127[214], stage127[215], stage127[216], stage127[217]},
      {stage129[39], stage128[52], stage127[259], stage126[248], stage125[259]}
   );
   gpc606_5 gpc606_5_7321(
      {stage125[223], stage125[224], stage125[225], stage125[226], stage125[227], stage125[228]},
      {stage127[218], stage127[219], stage127[220], stage127[221], stage127[222], stage127[223]},
      {stage129[40], stage128[53], stage127[260], stage126[249], stage125[260]}
   );
   gpc606_5 gpc606_5_7322(
      {stage125[229], stage125[230], stage125[231], stage125[232], stage125[233], stage125[234]},
      {stage127[224], stage127[225], stage127[226], stage127[227], stage127[228], stage127[229]},
      {stage129[41], stage128[54], stage127[261], stage126[250], stage125[261]}
   );
   gpc606_5 gpc606_5_7323(
      {stage125[235], stage125[236], stage125[237], stage125[238], stage125[239], stage125[240]},
      {stage127[230], stage127[231], stage127[232], stage127[233], stage127[234], stage127[235]},
      {stage129[42], stage128[55], stage127[262], stage126[251], stage125[262]}
   );
   gpc1_1 gpc1_1_7324(
      {stage126[219]},
      {stage126[252]}
   );
   gpc1_1 gpc1_1_7325(
      {stage126[220]},
      {stage126[253]}
   );
   gpc1_1 gpc1_1_7326(
      {stage126[221]},
      {stage126[254]}
   );
   gpc1_1 gpc1_1_7327(
      {stage126[222]},
      {stage126[255]}
   );
   gpc1_1 gpc1_1_7328(
      {stage126[223]},
      {stage126[256]}
   );
   gpc1_1 gpc1_1_7329(
      {stage126[224]},
      {stage126[257]}
   );
   gpc1_1 gpc1_1_7330(
      {stage126[225]},
      {stage126[258]}
   );
   gpc1_1 gpc1_1_7331(
      {stage126[226]},
      {stage126[259]}
   );
   gpc1_1 gpc1_1_7332(
      {stage126[227]},
      {stage126[260]}
   );
   gpc7_3 gpc7_3_7333(
      {stage126[228], stage126[229], stage126[230], stage126[231], stage126[232], stage126[233], stage126[234]},
      {stage128[56], stage127[263], stage126[261]}
   );
   gpc7_3 gpc7_3_7334(
      {stage126[235], stage126[236], stage126[237], stage126[238], stage126[239], stage126[240], stage126[241]},
      {stage128[57], stage127[264], stage126[262]}
   );
   gpc606_5 gpc606_5_7335(
      {stage127[236], stage127[237], stage127[238], stage127[239], stage127[240], stage127[241]},
      {stage129[12], stage129[13], stage129[14], stage129[15], stage129[16], stage129[17]},
      {stage131[0], stage130[5], stage129[43], stage128[58], stage127[265]}
   );
   gpc606_5 gpc606_5_7336(
      {stage127[242], stage127[243], stage127[244], stage127[245], stage127[246], stage127[247]},
      {stage129[18], stage129[19], stage129[20], stage129[21], stage129[22], stage129[23]},
      {stage131[1], stage130[6], stage129[44], stage128[59], stage127[266]}
   );
   gpc606_5 gpc606_5_7337(
      {stage127[248], stage127[249], stage127[250], stage127[251], stage127[252], stage127[253]},
      {stage129[24], stage129[25], stage129[26], stage129[27], stage129[28], stage129[29]},
      {stage131[2], stage130[7], stage129[45], stage128[60], stage127[267]}
   );
   gpc1_1 gpc1_1_7338(
      {stage128[31]},
      {stage128[61]}
   );
   gpc1_1 gpc1_1_7339(
      {stage128[32]},
      {stage128[62]}
   );
   gpc1_1 gpc1_1_7340(
      {stage128[33]},
      {stage128[63]}
   );
   gpc1_1 gpc1_1_7341(
      {stage128[34]},
      {stage128[64]}
   );
   gpc1_1 gpc1_1_7342(
      {stage128[35]},
      {stage128[65]}
   );
   gpc1_1 gpc1_1_7343(
      {stage128[36]},
      {stage128[66]}
   );
   gpc1_1 gpc1_1_7344(
      {stage128[37]},
      {stage128[67]}
   );
   gpc1_1 gpc1_1_7345(
      {stage128[38]},
      {stage128[68]}
   );
   gpc1_1 gpc1_1_7346(
      {stage128[39]},
      {stage128[69]}
   );
   gpc1_1 gpc1_1_7347(
      {stage128[40]},
      {stage128[70]}
   );
   gpc606_5 gpc606_5_7348(
      {stage128[41], stage128[42], stage128[43], stage128[44], stage128[45], stage128[46]},
      {stage130[0], stage130[1], stage130[2], stage130[3], stage130[4], 1'h0},
      {stage132[0], stage131[3], stage130[8], stage129[46], stage128[71]}
   );
   gpc1_1 gpc1_1_7349(
      {stage129[30]},
      {stage129[47]}
   );
   gpc1_1 gpc1_1_7350(
      {stage129[31]},
      {stage129[48]}
   );
   gpc1_1 gpc1_1_7351(
      {stage129[32]},
      {stage129[49]}
   );
   gpc1_1 gpc1_1_7352(
      {stage129[33]},
      {stage129[50]}
   );
   gpc1_1 gpc1_1_7353(
      {stage129[34]},
      {stage129[51]}
   );
   gpc1_1 gpc1_1_7354(
      {stage129[35]},
      {stage129[52]}
   );
   gpc1_1 gpc1_1_7355(
      {stage129[36]},
      {stage129[53]}
   );
   gpc1_1 gpc1_1_7356(
      {stage129[37]},
      {stage129[54]}
   );
   gpc1_1 gpc1_1_7357(
      {stage129[38]},
      {stage129[55]}
   );
   gpc1_1 gpc1_1_7358(
      {stage000[180]},
      {stage000[186]}
   );
   gpc615_5 gpc615_5_7359(
      {stage000[181], stage000[182], stage000[183], stage000[184], stage000[185]},
      {stage001[210]},
      {stage002[219], stage002[220], stage002[221], stage002[222], stage002[223], stage002[224]},
      {stage004[252], stage003[206], stage002[235], stage001[218], stage000[187]}
   );
   gpc1_1 gpc1_1_7360(
      {stage001[211]},
      {stage001[219]}
   );
   gpc1_1 gpc1_1_7361(
      {stage001[212]},
      {stage001[220]}
   );
   gpc1_1 gpc1_1_7362(
      {stage001[213]},
      {stage001[221]}
   );
   gpc1_1 gpc1_1_7363(
      {stage001[214]},
      {stage001[222]}
   );
   gpc1_1 gpc1_1_7364(
      {stage001[215]},
      {stage001[223]}
   );
   gpc1_1 gpc1_1_7365(
      {stage001[216]},
      {stage001[224]}
   );
   gpc1_1 gpc1_1_7366(
      {stage001[217]},
      {stage001[225]}
   );
   gpc1_1 gpc1_1_7367(
      {stage002[225]},
      {stage002[236]}
   );
   gpc1_1 gpc1_1_7368(
      {stage002[226]},
      {stage002[237]}
   );
   gpc1_1 gpc1_1_7369(
      {stage002[227]},
      {stage002[238]}
   );
   gpc1_1 gpc1_1_7370(
      {stage002[228]},
      {stage002[239]}
   );
   gpc1_1 gpc1_1_7371(
      {stage002[229]},
      {stage002[240]}
   );
   gpc2135_5 gpc2135_5_7372(
      {stage002[230], stage002[231], stage002[232], stage002[233], stage002[234]},
      {stage003[197], stage003[198], stage003[199]},
      {stage004[232]},
      {stage005[245], stage005[246]},
      {stage006[245], stage005[263], stage004[253], stage003[207], stage002[241]}
   );
   gpc1_1 gpc1_1_7373(
      {stage003[200]},
      {stage003[208]}
   );
   gpc1_1 gpc1_1_7374(
      {stage003[201]},
      {stage003[209]}
   );
   gpc1_1 gpc1_1_7375(
      {stage003[202]},
      {stage003[210]}
   );
   gpc1_1 gpc1_1_7376(
      {stage003[203]},
      {stage003[211]}
   );
   gpc1_1 gpc1_1_7377(
      {stage003[204]},
      {stage003[212]}
   );
   gpc1_1 gpc1_1_7378(
      {stage003[205]},
      {stage003[213]}
   );
   gpc1_1 gpc1_1_7379(
      {stage004[233]},
      {stage004[254]}
   );
   gpc1_1 gpc1_1_7380(
      {stage004[234]},
      {stage004[255]}
   );
   gpc1_1 gpc1_1_7381(
      {stage004[235]},
      {stage004[256]}
   );
   gpc1_1 gpc1_1_7382(
      {stage004[236]},
      {stage004[257]}
   );
   gpc1_1 gpc1_1_7383(
      {stage004[237]},
      {stage004[258]}
   );
   gpc1_1 gpc1_1_7384(
      {stage004[238]},
      {stage004[259]}
   );
   gpc1_1 gpc1_1_7385(
      {stage004[239]},
      {stage004[260]}
   );
   gpc606_5 gpc606_5_7386(
      {stage004[240], stage004[241], stage004[242], stage004[243], stage004[244], stage004[245]},
      {stage006[226], stage006[227], stage006[228], stage006[229], stage006[230], stage006[231]},
      {stage008[223], stage007[244], stage006[246], stage005[264], stage004[261]}
   );
   gpc606_5 gpc606_5_7387(
      {stage004[246], stage004[247], stage004[248], stage004[249], stage004[250], stage004[251]},
      {stage006[232], stage006[233], stage006[234], stage006[235], stage006[236], stage006[237]},
      {stage008[224], stage007[245], stage006[247], stage005[265], stage004[262]}
   );
   gpc1_1 gpc1_1_7388(
      {stage005[247]},
      {stage005[266]}
   );
   gpc1_1 gpc1_1_7389(
      {stage005[248]},
      {stage005[267]}
   );
   gpc1_1 gpc1_1_7390(
      {stage005[249]},
      {stage005[268]}
   );
   gpc1_1 gpc1_1_7391(
      {stage005[250]},
      {stage005[269]}
   );
   gpc1_1 gpc1_1_7392(
      {stage005[251]},
      {stage005[270]}
   );
   gpc1_1 gpc1_1_7393(
      {stage005[252]},
      {stage005[271]}
   );
   gpc1_1 gpc1_1_7394(
      {stage005[253]},
      {stage005[272]}
   );
   gpc1_1 gpc1_1_7395(
      {stage005[254]},
      {stage005[273]}
   );
   gpc1_1 gpc1_1_7396(
      {stage005[255]},
      {stage005[274]}
   );
   gpc1_1 gpc1_1_7397(
      {stage005[256]},
      {stage005[275]}
   );
   gpc606_5 gpc606_5_7398(
      {stage005[257], stage005[258], stage005[259], stage005[260], stage005[261], stage005[262]},
      {stage007[228], stage007[229], stage007[230], stage007[231], stage007[232], stage007[233]},
      {stage009[231], stage008[225], stage007[246], stage006[248], stage005[276]}
   );
   gpc1_1 gpc1_1_7399(
      {stage006[238]},
      {stage006[249]}
   );
   gpc606_5 gpc606_5_7400(
      {stage006[239], stage006[240], stage006[241], stage006[242], stage006[243], stage006[244]},
      {stage008[205], stage008[206], stage008[207], stage008[208], stage008[209], stage008[210]},
      {stage010[279], stage009[232], stage008[226], stage007[247], stage006[250]}
   );
   gpc606_5 gpc606_5_7401(
      {stage007[234], stage007[235], stage007[236], stage007[237], stage007[238], stage007[239]},
      {stage009[213], stage009[214], stage009[215], stage009[216], stage009[217], stage009[218]},
      {stage011[239], stage010[280], stage009[233], stage008[227], stage007[248]}
   );
   gpc615_5 gpc615_5_7402(
      {stage007[240], stage007[241], stage007[242], stage007[243], 1'h0},
      {stage008[211]},
      {stage009[219], stage009[220], stage009[221], stage009[222], stage009[223], stage009[224]},
      {stage011[240], stage010[281], stage009[234], stage008[228], stage007[249]}
   );
   gpc1_1 gpc1_1_7403(
      {stage008[212]},
      {stage008[229]}
   );
   gpc1_1 gpc1_1_7404(
      {stage008[213]},
      {stage008[230]}
   );
   gpc1_1 gpc1_1_7405(
      {stage008[214]},
      {stage008[231]}
   );
   gpc1_1 gpc1_1_7406(
      {stage008[215]},
      {stage008[232]}
   );
   gpc1_1 gpc1_1_7407(
      {stage008[216]},
      {stage008[233]}
   );
   gpc1_1 gpc1_1_7408(
      {stage008[217]},
      {stage008[234]}
   );
   gpc615_5 gpc615_5_7409(
      {stage008[218], stage008[219], stage008[220], stage008[221], stage008[222]},
      {stage009[225]},
      {stage010[257], stage010[258], stage010[259], stage010[260], stage010[261], stage010[262]},
      {stage012[310], stage011[241], stage010[282], stage009[235], stage008[235]}
   );
   gpc615_5 gpc615_5_7410(
      {stage009[226], stage009[227], stage009[228], stage009[229], stage009[230]},
      {stage010[263]},
      {stage011[220], stage011[221], stage011[222], stage011[223], stage011[224], stage011[225]},
      {stage013[235], stage012[311], stage011[242], stage010[283], stage009[236]}
   );
   gpc1_1 gpc1_1_7411(
      {stage010[264]},
      {stage010[284]}
   );
   gpc1_1 gpc1_1_7412(
      {stage010[265]},
      {stage010[285]}
   );
   gpc1_1 gpc1_1_7413(
      {stage010[266]},
      {stage010[286]}
   );
   gpc1_1 gpc1_1_7414(
      {stage010[267]},
      {stage010[287]}
   );
   gpc1_1 gpc1_1_7415(
      {stage010[268]},
      {stage010[288]}
   );
   gpc615_5 gpc615_5_7416(
      {stage010[269], stage010[270], stage010[271], stage010[272], stage010[273]},
      {stage011[226]},
      {stage012[277], stage012[278], stage012[279], stage012[280], stage012[281], stage012[282]},
      {stage014[288], stage013[236], stage012[312], stage011[243], stage010[289]}
   );
   gpc615_5 gpc615_5_7417(
      {stage010[274], stage010[275], stage010[276], stage010[277], stage010[278]},
      {stage011[227]},
      {stage012[283], stage012[284], stage012[285], stage012[286], stage012[287], stage012[288]},
      {stage014[289], stage013[237], stage012[313], stage011[244], stage010[290]}
   );
   gpc1_1 gpc1_1_7418(
      {stage011[228]},
      {stage011[245]}
   );
   gpc1_1 gpc1_1_7419(
      {stage011[229]},
      {stage011[246]}
   );
   gpc1_1 gpc1_1_7420(
      {stage011[230]},
      {stage011[247]}
   );
   gpc1_1 gpc1_1_7421(
      {stage011[231]},
      {stage011[248]}
   );
   gpc1_1 gpc1_1_7422(
      {stage011[232]},
      {stage011[249]}
   );
   gpc1_1 gpc1_1_7423(
      {stage011[233]},
      {stage011[250]}
   );
   gpc1_1 gpc1_1_7424(
      {stage011[234]},
      {stage011[251]}
   );
   gpc1_1 gpc1_1_7425(
      {stage011[235]},
      {stage011[252]}
   );
   gpc623_5 gpc623_5_7426(
      {stage011[236], stage011[237], stage011[238]},
      {stage012[289], stage012[290]},
      {stage013[208], stage013[209], stage013[210], stage013[211], stage013[212], stage013[213]},
      {stage015[240], stage014[290], stage013[238], stage012[314], stage011[253]}
   );
   gpc1_1 gpc1_1_7427(
      {stage012[291]},
      {stage012[315]}
   );
   gpc606_5 gpc606_5_7428(
      {stage012[292], stage012[293], stage012[294], stage012[295], stage012[296], stage012[297]},
      {stage014[258], stage014[259], stage014[260], stage014[261], stage014[262], stage014[263]},
      {stage016[275], stage015[241], stage014[291], stage013[239], stage012[316]}
   );
   gpc606_5 gpc606_5_7429(
      {stage012[298], stage012[299], stage012[300], stage012[301], stage012[302], stage012[303]},
      {stage014[264], stage014[265], stage014[266], stage014[267], stage014[268], stage014[269]},
      {stage016[276], stage015[242], stage014[292], stage013[240], stage012[317]}
   );
   gpc606_5 gpc606_5_7430(
      {stage012[304], stage012[305], stage012[306], stage012[307], stage012[308], stage012[309]},
      {stage014[270], stage014[271], stage014[272], stage014[273], stage014[274], stage014[275]},
      {stage016[277], stage015[243], stage014[293], stage013[241], stage012[318]}
   );
   gpc1_1 gpc1_1_7431(
      {stage013[214]},
      {stage013[242]}
   );
   gpc1_1 gpc1_1_7432(
      {stage013[215]},
      {stage013[243]}
   );
   gpc1_1 gpc1_1_7433(
      {stage013[216]},
      {stage013[244]}
   );
   gpc1_1 gpc1_1_7434(
      {stage013[217]},
      {stage013[245]}
   );
   gpc1_1 gpc1_1_7435(
      {stage013[218]},
      {stage013[246]}
   );
   gpc1_1 gpc1_1_7436(
      {stage013[219]},
      {stage013[247]}
   );
   gpc1_1 gpc1_1_7437(
      {stage013[220]},
      {stage013[248]}
   );
   gpc1_1 gpc1_1_7438(
      {stage013[221]},
      {stage013[249]}
   );
   gpc1_1 gpc1_1_7439(
      {stage013[222]},
      {stage013[250]}
   );
   gpc606_5 gpc606_5_7440(
      {stage013[223], stage013[224], stage013[225], stage013[226], stage013[227], stage013[228]},
      {stage015[223], stage015[224], stage015[225], stage015[226], stage015[227], stage015[228]},
      {stage017[266], stage016[278], stage015[244], stage014[294], stage013[251]}
   );
   gpc606_5 gpc606_5_7441(
      {stage013[229], stage013[230], stage013[231], stage013[232], stage013[233], stage013[234]},
      {stage015[229], stage015[230], stage015[231], stage015[232], stage015[233], stage015[234]},
      {stage017[267], stage016[279], stage015[245], stage014[295], stage013[252]}
   );
   gpc606_5 gpc606_5_7442(
      {stage014[276], stage014[277], stage014[278], stage014[279], stage014[280], stage014[281]},
      {stage016[246], stage016[247], stage016[248], stage016[249], stage016[250], stage016[251]},
      {stage018[241], stage017[268], stage016[280], stage015[246], stage014[296]}
   );
   gpc606_5 gpc606_5_7443(
      {stage014[282], stage014[283], stage014[284], stage014[285], stage014[286], stage014[287]},
      {stage016[252], stage016[253], stage016[254], stage016[255], stage016[256], stage016[257]},
      {stage018[242], stage017[269], stage016[281], stage015[247], stage014[297]}
   );
   gpc1_1 gpc1_1_7444(
      {stage015[235]},
      {stage015[248]}
   );
   gpc1_1 gpc1_1_7445(
      {stage015[236]},
      {stage015[249]}
   );
   gpc1_1 gpc1_1_7446(
      {stage015[237]},
      {stage015[250]}
   );
   gpc1_1 gpc1_1_7447(
      {stage015[238]},
      {stage015[251]}
   );
   gpc1_1 gpc1_1_7448(
      {stage015[239]},
      {stage015[252]}
   );
   gpc606_5 gpc606_5_7449(
      {stage016[258], stage016[259], stage016[260], stage016[261], stage016[262], stage016[263]},
      {stage018[222], stage018[223], stage018[224], stage018[225], stage018[226], stage018[227]},
      {stage020[219], stage019[246], stage018[243], stage017[270], stage016[282]}
   );
   gpc606_5 gpc606_5_7450(
      {stage016[264], stage016[265], stage016[266], stage016[267], stage016[268], stage016[269]},
      {stage018[228], stage018[229], stage018[230], stage018[231], stage018[232], stage018[233]},
      {stage020[220], stage019[247], stage018[244], stage017[271], stage016[283]}
   );
   gpc606_5 gpc606_5_7451(
      {stage016[270], stage016[271], stage016[272], stage016[273], stage016[274], 1'h0},
      {stage018[234], stage018[235], stage018[236], stage018[237], stage018[238], stage018[239]},
      {stage020[221], stage019[248], stage018[245], stage017[272], stage016[284]}
   );
   gpc1_1 gpc1_1_7452(
      {stage017[251]},
      {stage017[273]}
   );
   gpc1_1 gpc1_1_7453(
      {stage017[252]},
      {stage017[274]}
   );
   gpc1_1 gpc1_1_7454(
      {stage017[253]},
      {stage017[275]}
   );
   gpc606_5 gpc606_5_7455(
      {stage017[254], stage017[255], stage017[256], stage017[257], stage017[258], stage017[259]},
      {stage019[222], stage019[223], stage019[224], stage019[225], stage019[226], stage019[227]},
      {stage021[271], stage020[222], stage019[249], stage018[246], stage017[276]}
   );
   gpc606_5 gpc606_5_7456(
      {stage017[260], stage017[261], stage017[262], stage017[263], stage017[264], stage017[265]},
      {stage019[228], stage019[229], stage019[230], stage019[231], stage019[232], stage019[233]},
      {stage021[272], stage020[223], stage019[250], stage018[247], stage017[277]}
   );
   gpc1_1 gpc1_1_7457(
      {stage018[240]},
      {stage018[248]}
   );
   gpc1_1 gpc1_1_7458(
      {stage019[234]},
      {stage019[251]}
   );
   gpc1_1 gpc1_1_7459(
      {stage019[235]},
      {stage019[252]}
   );
   gpc1_1 gpc1_1_7460(
      {stage019[236]},
      {stage019[253]}
   );
   gpc1_1 gpc1_1_7461(
      {stage019[237]},
      {stage019[254]}
   );
   gpc1_1 gpc1_1_7462(
      {stage019[238]},
      {stage019[255]}
   );
   gpc1_1 gpc1_1_7463(
      {stage019[239]},
      {stage019[256]}
   );
   gpc606_5 gpc606_5_7464(
      {stage019[240], stage019[241], stage019[242], stage019[243], stage019[244], stage019[245]},
      {stage021[239], stage021[240], stage021[241], stage021[242], stage021[243], stage021[244]},
      {stage023[295], stage022[215], stage021[273], stage020[224], stage019[257]}
   );
   gpc1_1 gpc1_1_7465(
      {stage020[211]},
      {stage020[225]}
   );
   gpc1_1 gpc1_1_7466(
      {stage020[212]},
      {stage020[226]}
   );
   gpc1_1 gpc1_1_7467(
      {stage020[213]},
      {stage020[227]}
   );
   gpc1325_5 gpc1325_5_7468(
      {stage020[214], stage020[215], stage020[216], stage020[217], stage020[218]},
      {stage021[245], stage021[246]},
      {stage022[201], stage022[202], stage022[203]},
      {stage023[265]},
      {stage024[245], stage023[296], stage022[216], stage021[274], stage020[228]}
   );
   gpc1_1 gpc1_1_7469(
      {stage021[247]},
      {stage021[275]}
   );
   gpc1_1 gpc1_1_7470(
      {stage021[248]},
      {stage021[276]}
   );
   gpc1_1 gpc1_1_7471(
      {stage021[249]},
      {stage021[277]}
   );
   gpc1_1 gpc1_1_7472(
      {stage021[250]},
      {stage021[278]}
   );
   gpc1_1 gpc1_1_7473(
      {stage021[251]},
      {stage021[279]}
   );
   gpc1_1 gpc1_1_7474(
      {stage021[252]},
      {stage021[280]}
   );
   gpc1_1 gpc1_1_7475(
      {stage021[253]},
      {stage021[281]}
   );
   gpc606_5 gpc606_5_7476(
      {stage021[254], stage021[255], stage021[256], stage021[257], stage021[258], stage021[259]},
      {stage023[266], stage023[267], stage023[268], stage023[269], stage023[270], stage023[271]},
      {stage025[279], stage024[246], stage023[297], stage022[217], stage021[282]}
   );
   gpc606_5 gpc606_5_7477(
      {stage021[260], stage021[261], stage021[262], stage021[263], stage021[264], stage021[265]},
      {stage023[272], stage023[273], stage023[274], stage023[275], stage023[276], stage023[277]},
      {stage025[280], stage024[247], stage023[298], stage022[218], stage021[283]}
   );
   gpc1415_5 gpc1415_5_7478(
      {stage021[266], stage021[267], stage021[268], stage021[269], stage021[270]},
      {stage022[204]},
      {stage023[278], stage023[279], stage023[280], stage023[281]},
      {stage024[225]},
      {stage025[281], stage024[248], stage023[299], stage022[219], stage021[284]}
   );
   gpc1_1 gpc1_1_7479(
      {stage022[205]},
      {stage022[220]}
   );
   gpc1_1 gpc1_1_7480(
      {stage022[206]},
      {stage022[221]}
   );
   gpc1_1 gpc1_1_7481(
      {stage022[207]},
      {stage022[222]}
   );
   gpc1_1 gpc1_1_7482(
      {stage022[208]},
      {stage022[223]}
   );
   gpc606_5 gpc606_5_7483(
      {stage022[209], stage022[210], stage022[211], stage022[212], stage022[213], stage022[214]},
      {stage024[226], stage024[227], stage024[228], stage024[229], stage024[230], stage024[231]},
      {stage026[234], stage025[282], stage024[249], stage023[300], stage022[224]}
   );
   gpc1_1 gpc1_1_7484(
      {stage023[282]},
      {stage023[301]}
   );
   gpc1_1 gpc1_1_7485(
      {stage023[283]},
      {stage023[302]}
   );
   gpc1_1 gpc1_1_7486(
      {stage023[284]},
      {stage023[303]}
   );
   gpc1_1 gpc1_1_7487(
      {stage023[285]},
      {stage023[304]}
   );
   gpc1_1 gpc1_1_7488(
      {stage023[286]},
      {stage023[305]}
   );
   gpc1_1 gpc1_1_7489(
      {stage023[287]},
      {stage023[306]}
   );
   gpc1_1 gpc1_1_7490(
      {stage023[288]},
      {stage023[307]}
   );
   gpc606_5 gpc606_5_7491(
      {stage023[289], stage023[290], stage023[291], stage023[292], stage023[293], stage023[294]},
      {stage025[257], stage025[258], stage025[259], stage025[260], stage025[261], stage025[262]},
      {stage027[229], stage026[235], stage025[283], stage024[250], stage023[308]}
   );
   gpc1_1 gpc1_1_7492(
      {stage024[232]},
      {stage024[251]}
   );
   gpc606_5 gpc606_5_7493(
      {stage024[233], stage024[234], stage024[235], stage024[236], stage024[237], stage024[238]},
      {stage026[222], stage026[223], stage026[224], stage026[225], stage026[226], stage026[227]},
      {stage028[239], stage027[230], stage026[236], stage025[284], stage024[252]}
   );
   gpc606_5 gpc606_5_7494(
      {stage024[239], stage024[240], stage024[241], stage024[242], stage024[243], stage024[244]},
      {stage026[228], stage026[229], stage026[230], stage026[231], stage026[232], stage026[233]},
      {stage028[240], stage027[231], stage026[237], stage025[285], stage024[253]}
   );
   gpc1_1 gpc1_1_7495(
      {stage025[263]},
      {stage025[286]}
   );
   gpc1_1 gpc1_1_7496(
      {stage025[264]},
      {stage025[287]}
   );
   gpc1_1 gpc1_1_7497(
      {stage025[265]},
      {stage025[288]}
   );
   gpc1_1 gpc1_1_7498(
      {stage025[266]},
      {stage025[289]}
   );
   gpc606_5 gpc606_5_7499(
      {stage025[267], stage025[268], stage025[269], stage025[270], stage025[271], stage025[272]},
      {stage027[211], stage027[212], stage027[213], stage027[214], stage027[215], stage027[216]},
      {stage029[274], stage028[241], stage027[232], stage026[238], stage025[290]}
   );
   gpc606_5 gpc606_5_7500(
      {stage025[273], stage025[274], stage025[275], stage025[276], stage025[277], stage025[278]},
      {stage027[217], stage027[218], stage027[219], stage027[220], stage027[221], stage027[222]},
      {stage029[275], stage028[242], stage027[233], stage026[239], stage025[291]}
   );
   gpc606_5 gpc606_5_7501(
      {stage027[223], stage027[224], stage027[225], stage027[226], stage027[227], stage027[228]},
      {stage029[251], stage029[252], stage029[253], stage029[254], stage029[255], stage029[256]},
      {stage031[238], stage030[230], stage029[276], stage028[243], stage027[234]}
   );
   gpc1_1 gpc1_1_7502(
      {stage028[224]},
      {stage028[244]}
   );
   gpc1_1 gpc1_1_7503(
      {stage028[225]},
      {stage028[245]}
   );
   gpc1_1 gpc1_1_7504(
      {stage028[226]},
      {stage028[246]}
   );
   gpc1_1 gpc1_1_7505(
      {stage028[227]},
      {stage028[247]}
   );
   gpc1_1 gpc1_1_7506(
      {stage028[228]},
      {stage028[248]}
   );
   gpc1_1 gpc1_1_7507(
      {stage028[229]},
      {stage028[249]}
   );
   gpc1_1 gpc1_1_7508(
      {stage028[230]},
      {stage028[250]}
   );
   gpc1_1 gpc1_1_7509(
      {stage028[231]},
      {stage028[251]}
   );
   gpc1_1 gpc1_1_7510(
      {stage028[232]},
      {stage028[252]}
   );
   gpc606_5 gpc606_5_7511(
      {stage028[233], stage028[234], stage028[235], stage028[236], stage028[237], stage028[238]},
      {stage030[210], stage030[211], stage030[212], stage030[213], stage030[214], stage030[215]},
      {stage032[284], stage031[239], stage030[231], stage029[277], stage028[253]}
   );
   gpc1_1 gpc1_1_7512(
      {stage029[257]},
      {stage029[278]}
   );
   gpc1_1 gpc1_1_7513(
      {stage029[258]},
      {stage029[279]}
   );
   gpc1_1 gpc1_1_7514(
      {stage029[259]},
      {stage029[280]}
   );
   gpc1_1 gpc1_1_7515(
      {stage029[260]},
      {stage029[281]}
   );
   gpc1_1 gpc1_1_7516(
      {stage029[261]},
      {stage029[282]}
   );
   gpc606_5 gpc606_5_7517(
      {stage029[262], stage029[263], stage029[264], stage029[265], stage029[266], stage029[267]},
      {stage031[210], stage031[211], stage031[212], stage031[213], stage031[214], stage031[215]},
      {stage033[284], stage032[285], stage031[240], stage030[232], stage029[283]}
   );
   gpc606_5 gpc606_5_7518(
      {stage029[268], stage029[269], stage029[270], stage029[271], stage029[272], stage029[273]},
      {stage031[216], stage031[217], stage031[218], stage031[219], stage031[220], stage031[221]},
      {stage033[285], stage032[286], stage031[241], stage030[233], stage029[284]}
   );
   gpc1_1 gpc1_1_7519(
      {stage030[216]},
      {stage030[234]}
   );
   gpc1_1 gpc1_1_7520(
      {stage030[217]},
      {stage030[235]}
   );
   gpc1_1 gpc1_1_7521(
      {stage030[218]},
      {stage030[236]}
   );
   gpc1_1 gpc1_1_7522(
      {stage030[219]},
      {stage030[237]}
   );
   gpc615_5 gpc615_5_7523(
      {stage030[220], stage030[221], stage030[222], stage030[223], stage030[224]},
      {stage031[222]},
      {stage032[263], stage032[264], stage032[265], stage032[266], stage032[267], stage032[268]},
      {stage034[280], stage033[286], stage032[287], stage031[242], stage030[238]}
   );
   gpc615_5 gpc615_5_7524(
      {stage030[225], stage030[226], stage030[227], stage030[228], stage030[229]},
      {stage031[223]},
      {stage032[269], stage032[270], stage032[271], stage032[272], stage032[273], stage032[274]},
      {stage034[281], stage033[287], stage032[288], stage031[243], stage030[239]}
   );
   gpc1_1 gpc1_1_7525(
      {stage031[224]},
      {stage031[244]}
   );
   gpc1_1 gpc1_1_7526(
      {stage031[225]},
      {stage031[245]}
   );
   gpc1_1 gpc1_1_7527(
      {stage031[226]},
      {stage031[246]}
   );
   gpc1_1 gpc1_1_7528(
      {stage031[227]},
      {stage031[247]}
   );
   gpc615_5 gpc615_5_7529(
      {stage031[228], stage031[229], stage031[230], stage031[231], stage031[232]},
      {stage032[275]},
      {stage033[266], stage033[267], stage033[268], stage033[269], stage033[270], stage033[271]},
      {stage035[254], stage034[282], stage033[288], stage032[289], stage031[248]}
   );
   gpc615_5 gpc615_5_7530(
      {stage031[233], stage031[234], stage031[235], stage031[236], stage031[237]},
      {stage032[276]},
      {stage033[272], stage033[273], stage033[274], stage033[275], stage033[276], stage033[277]},
      {stage035[255], stage034[283], stage033[289], stage032[290], stage031[249]}
   );
   gpc1_1 gpc1_1_7531(
      {stage032[277]},
      {stage032[291]}
   );
   gpc1_1 gpc1_1_7532(
      {stage032[278]},
      {stage032[292]}
   );
   gpc1_1 gpc1_1_7533(
      {stage032[279]},
      {stage032[293]}
   );
   gpc1_1 gpc1_1_7534(
      {stage032[280]},
      {stage032[294]}
   );
   gpc1_1 gpc1_1_7535(
      {stage032[281]},
      {stage032[295]}
   );
   gpc1_1 gpc1_1_7536(
      {stage032[282]},
      {stage032[296]}
   );
   gpc1_1 gpc1_1_7537(
      {stage032[283]},
      {stage032[297]}
   );
   gpc606_5 gpc606_5_7538(
      {stage033[278], stage033[279], stage033[280], stage033[281], stage033[282], stage033[283]},
      {stage035[237], stage035[238], stage035[239], stage035[240], stage035[241], stage035[242]},
      {stage037[259], stage036[216], stage035[256], stage034[284], stage033[290]}
   );
   gpc1_1 gpc1_1_7539(
      {stage034[262]},
      {stage034[285]}
   );
   gpc1_1 gpc1_1_7540(
      {stage034[263]},
      {stage034[286]}
   );
   gpc1_1 gpc1_1_7541(
      {stage034[264]},
      {stage034[287]}
   );
   gpc1_1 gpc1_1_7542(
      {stage034[265]},
      {stage034[288]}
   );
   gpc1_1 gpc1_1_7543(
      {stage034[266]},
      {stage034[289]}
   );
   gpc1_1 gpc1_1_7544(
      {stage034[267]},
      {stage034[290]}
   );
   gpc1_1 gpc1_1_7545(
      {stage034[268]},
      {stage034[291]}
   );
   gpc1_1 gpc1_1_7546(
      {stage034[269]},
      {stage034[292]}
   );
   gpc1_1 gpc1_1_7547(
      {stage034[270]},
      {stage034[293]}
   );
   gpc1_1 gpc1_1_7548(
      {stage034[271]},
      {stage034[294]}
   );
   gpc1_1 gpc1_1_7549(
      {stage034[272]},
      {stage034[295]}
   );
   gpc1_1 gpc1_1_7550(
      {stage034[273]},
      {stage034[296]}
   );
   gpc1_1 gpc1_1_7551(
      {stage034[274]},
      {stage034[297]}
   );
   gpc615_5 gpc615_5_7552(
      {stage034[275], stage034[276], stage034[277], stage034[278], stage034[279]},
      {stage035[243]},
      {stage036[203], stage036[204], stage036[205], stage036[206], stage036[207], stage036[208]},
      {stage038[234], stage037[260], stage036[217], stage035[257], stage034[298]}
   );
   gpc615_5 gpc615_5_7553(
      {stage035[244], stage035[245], stage035[246], stage035[247], stage035[248]},
      {stage036[209]},
      {stage037[229], stage037[230], stage037[231], stage037[232], stage037[233], stage037[234]},
      {stage039[243], stage038[235], stage037[261], stage036[218], stage035[258]}
   );
   gpc615_5 gpc615_5_7554(
      {stage035[249], stage035[250], stage035[251], stage035[252], stage035[253]},
      {stage036[210]},
      {stage037[235], stage037[236], stage037[237], stage037[238], stage037[239], stage037[240]},
      {stage039[244], stage038[236], stage037[262], stage036[219], stage035[259]}
   );
   gpc1_1 gpc1_1_7555(
      {stage036[211]},
      {stage036[220]}
   );
   gpc1_1 gpc1_1_7556(
      {stage036[212]},
      {stage036[221]}
   );
   gpc1_1 gpc1_1_7557(
      {stage036[213]},
      {stage036[222]}
   );
   gpc1_1 gpc1_1_7558(
      {stage036[214]},
      {stage036[223]}
   );
   gpc1_1 gpc1_1_7559(
      {stage036[215]},
      {stage036[224]}
   );
   gpc1_1 gpc1_1_7560(
      {stage037[241]},
      {stage037[263]}
   );
   gpc1_1 gpc1_1_7561(
      {stage037[242]},
      {stage037[264]}
   );
   gpc1_1 gpc1_1_7562(
      {stage037[243]},
      {stage037[265]}
   );
   gpc1_1 gpc1_1_7563(
      {stage037[244]},
      {stage037[266]}
   );
   gpc1_1 gpc1_1_7564(
      {stage037[245]},
      {stage037[267]}
   );
   gpc1_1 gpc1_1_7565(
      {stage037[246]},
      {stage037[268]}
   );
   gpc606_5 gpc606_5_7566(
      {stage037[247], stage037[248], stage037[249], stage037[250], stage037[251], stage037[252]},
      {stage039[224], stage039[225], stage039[226], stage039[227], stage039[228], stage039[229]},
      {stage041[253], stage040[286], stage039[245], stage038[237], stage037[269]}
   );
   gpc606_5 gpc606_5_7567(
      {stage037[253], stage037[254], stage037[255], stage037[256], stage037[257], stage037[258]},
      {stage039[230], stage039[231], stage039[232], stage039[233], stage039[234], stage039[235]},
      {stage041[254], stage040[287], stage039[246], stage038[238], stage037[270]}
   );
   gpc1_1 gpc1_1_7568(
      {stage038[223]},
      {stage038[239]}
   );
   gpc1_1 gpc1_1_7569(
      {stage038[224]},
      {stage038[240]}
   );
   gpc1_1 gpc1_1_7570(
      {stage038[225]},
      {stage038[241]}
   );
   gpc1_1 gpc1_1_7571(
      {stage038[226]},
      {stage038[242]}
   );
   gpc1_1 gpc1_1_7572(
      {stage038[227]},
      {stage038[243]}
   );
   gpc1_1 gpc1_1_7573(
      {stage038[228]},
      {stage038[244]}
   );
   gpc1_1 gpc1_1_7574(
      {stage038[229]},
      {stage038[245]}
   );
   gpc1_1 gpc1_1_7575(
      {stage038[230]},
      {stage038[246]}
   );
   gpc1_1 gpc1_1_7576(
      {stage038[231]},
      {stage038[247]}
   );
   gpc1_1 gpc1_1_7577(
      {stage038[232]},
      {stage038[248]}
   );
   gpc1_1 gpc1_1_7578(
      {stage038[233]},
      {stage038[249]}
   );
   gpc1_1 gpc1_1_7579(
      {stage039[236]},
      {stage039[247]}
   );
   gpc1_1 gpc1_1_7580(
      {stage039[237]},
      {stage039[248]}
   );
   gpc615_5 gpc615_5_7581(
      {stage039[238], stage039[239], stage039[240], stage039[241], stage039[242]},
      {stage040[268]},
      {stage041[237], stage041[238], stage041[239], stage041[240], stage041[241], stage041[242]},
      {stage043[210], stage042[279], stage041[255], stage040[288], stage039[249]}
   );
   gpc1_1 gpc1_1_7582(
      {stage040[269]},
      {stage040[289]}
   );
   gpc1_1 gpc1_1_7583(
      {stage040[270]},
      {stage040[290]}
   );
   gpc1_1 gpc1_1_7584(
      {stage040[271]},
      {stage040[291]}
   );
   gpc1_1 gpc1_1_7585(
      {stage040[272]},
      {stage040[292]}
   );
   gpc1_1 gpc1_1_7586(
      {stage040[273]},
      {stage040[293]}
   );
   gpc1_1 gpc1_1_7587(
      {stage040[274]},
      {stage040[294]}
   );
   gpc1_1 gpc1_1_7588(
      {stage040[275]},
      {stage040[295]}
   );
   gpc1_1 gpc1_1_7589(
      {stage040[276]},
      {stage040[296]}
   );
   gpc1_1 gpc1_1_7590(
      {stage040[277]},
      {stage040[297]}
   );
   gpc1_1 gpc1_1_7591(
      {stage040[278]},
      {stage040[298]}
   );
   gpc1_1 gpc1_1_7592(
      {stage040[279]},
      {stage040[299]}
   );
   gpc606_5 gpc606_5_7593(
      {stage040[280], stage040[281], stage040[282], stage040[283], stage040[284], stage040[285]},
      {stage042[247], stage042[248], stage042[249], stage042[250], stage042[251], stage042[252]},
      {stage044[220], stage043[211], stage042[280], stage041[256], stage040[300]}
   );
   gpc1_1 gpc1_1_7594(
      {stage041[243]},
      {stage041[257]}
   );
   gpc1_1 gpc1_1_7595(
      {stage041[244]},
      {stage041[258]}
   );
   gpc1_1 gpc1_1_7596(
      {stage041[245]},
      {stage041[259]}
   );
   gpc1_1 gpc1_1_7597(
      {stage041[246]},
      {stage041[260]}
   );
   gpc1_1 gpc1_1_7598(
      {stage041[247]},
      {stage041[261]}
   );
   gpc1_1 gpc1_1_7599(
      {stage041[248]},
      {stage041[262]}
   );
   gpc1_1 gpc1_1_7600(
      {stage041[249]},
      {stage041[263]}
   );
   gpc1_1 gpc1_1_7601(
      {stage041[250]},
      {stage041[264]}
   );
   gpc1_1 gpc1_1_7602(
      {stage041[251]},
      {stage041[265]}
   );
   gpc1_1 gpc1_1_7603(
      {stage041[252]},
      {stage041[266]}
   );
   gpc1_1 gpc1_1_7604(
      {stage042[253]},
      {stage042[281]}
   );
   gpc1_1 gpc1_1_7605(
      {stage042[254]},
      {stage042[282]}
   );
   gpc1_1 gpc1_1_7606(
      {stage042[255]},
      {stage042[283]}
   );
   gpc1_1 gpc1_1_7607(
      {stage042[256]},
      {stage042[284]}
   );
   gpc1_1 gpc1_1_7608(
      {stage042[257]},
      {stage042[285]}
   );
   gpc1_1 gpc1_1_7609(
      {stage042[258]},
      {stage042[286]}
   );
   gpc1325_5 gpc1325_5_7610(
      {stage042[259], stage042[260], stage042[261], stage042[262], stage042[263]},
      {stage043[196], stage043[197]},
      {stage044[208], stage044[209], stage044[210]},
      {stage045[250]},
      {stage046[263], stage045[266], stage044[221], stage043[212], stage042[287]}
   );
   gpc1325_5 gpc1325_5_7611(
      {stage042[264], stage042[265], stage042[266], stage042[267], stage042[268]},
      {stage043[198], stage043[199]},
      {stage044[211], stage044[212], stage044[213]},
      {stage045[251]},
      {stage046[264], stage045[267], stage044[222], stage043[213], stage042[288]}
   );
   gpc1325_5 gpc1325_5_7612(
      {stage042[269], stage042[270], stage042[271], stage042[272], stage042[273]},
      {stage043[200], stage043[201]},
      {stage044[214], stage044[215], stage044[216]},
      {stage045[252]},
      {stage046[265], stage045[268], stage044[223], stage043[214], stage042[289]}
   );
   gpc1325_5 gpc1325_5_7613(
      {stage042[274], stage042[275], stage042[276], stage042[277], stage042[278]},
      {stage043[202], stage043[203]},
      {stage044[217], stage044[218], stage044[219]},
      {stage045[253]},
      {stage046[266], stage045[269], stage044[224], stage043[215], stage042[290]}
   );
   gpc606_5 gpc606_5_7614(
      {stage043[204], stage043[205], stage043[206], stage043[207], stage043[208], stage043[209]},
      {stage045[254], stage045[255], stage045[256], stage045[257], stage045[258], stage045[259]},
      {stage047[224], stage046[267], stage045[270], stage044[225], stage043[216]}
   );
   gpc606_5 gpc606_5_7615(
      {stage045[260], stage045[261], stage045[262], stage045[263], stage045[264], stage045[265]},
      {stage047[198], stage047[199], stage047[200], stage047[201], stage047[202], stage047[203]},
      {stage049[245], stage048[321], stage047[225], stage046[268], stage045[271]}
   );
   gpc615_5 gpc615_5_7616(
      {stage046[249], stage046[250], stage046[251], stage046[252], stage046[253]},
      {stage047[204]},
      {stage048[295], stage048[296], stage048[297], stage048[298], stage048[299], stage048[300]},
      {stage050[268], stage049[246], stage048[322], stage047[226], stage046[269]}
   );
   gpc615_5 gpc615_5_7617(
      {stage046[254], stage046[255], stage046[256], stage046[257], stage046[258]},
      {stage047[205]},
      {stage048[301], stage048[302], stage048[303], stage048[304], stage048[305], stage048[306]},
      {stage050[269], stage049[247], stage048[323], stage047[227], stage046[270]}
   );
   gpc615_5 gpc615_5_7618(
      {stage046[259], stage046[260], stage046[261], stage046[262], 1'h0},
      {stage047[206]},
      {stage048[307], stage048[308], stage048[309], stage048[310], stage048[311], stage048[312]},
      {stage050[270], stage049[248], stage048[324], stage047[228], stage046[271]}
   );
   gpc7_3 gpc7_3_7619(
      {stage047[207], stage047[208], stage047[209], stage047[210], stage047[211], stage047[212], stage047[213]},
      {stage049[249], stage048[325], stage047[229]}
   );
   gpc606_5 gpc606_5_7620(
      {stage047[214], stage047[215], stage047[216], stage047[217], stage047[218], stage047[219]},
      {stage049[230], stage049[231], stage049[232], stage049[233], stage049[234], stage049[235]},
      {stage051[237], stage050[271], stage049[250], stage048[326], stage047[230]}
   );
   gpc606_5 gpc606_5_7621(
      {stage047[220], stage047[221], stage047[222], stage047[223], 1'h0, 1'h0},
      {stage049[236], stage049[237], stage049[238], stage049[239], stage049[240], stage049[241]},
      {stage051[238], stage050[272], stage049[251], stage048[327], stage047[231]}
   );
   gpc1_1 gpc1_1_7622(
      {stage048[313]},
      {stage048[328]}
   );
   gpc1_1 gpc1_1_7623(
      {stage048[314]},
      {stage048[329]}
   );
   gpc1_1 gpc1_1_7624(
      {stage048[315]},
      {stage048[330]}
   );
   gpc1_1 gpc1_1_7625(
      {stage048[316]},
      {stage048[331]}
   );
   gpc1_1 gpc1_1_7626(
      {stage048[317]},
      {stage048[332]}
   );
   gpc1_1 gpc1_1_7627(
      {stage048[318]},
      {stage048[333]}
   );
   gpc1_1 gpc1_1_7628(
      {stage048[319]},
      {stage048[334]}
   );
   gpc1_1 gpc1_1_7629(
      {stage048[320]},
      {stage048[335]}
   );
   gpc1_1 gpc1_1_7630(
      {stage049[242]},
      {stage049[252]}
   );
   gpc1_1 gpc1_1_7631(
      {stage049[243]},
      {stage049[253]}
   );
   gpc1_1 gpc1_1_7632(
      {stage049[244]},
      {stage049[254]}
   );
   gpc1_1 gpc1_1_7633(
      {stage050[255]},
      {stage050[273]}
   );
   gpc1_1 gpc1_1_7634(
      {stage050[256]},
      {stage050[274]}
   );
   gpc1_1 gpc1_1_7635(
      {stage050[257]},
      {stage050[275]}
   );
   gpc615_5 gpc615_5_7636(
      {stage050[258], stage050[259], stage050[260], stage050[261], stage050[262]},
      {stage051[222]},
      {stage052[243], stage052[244], stage052[245], stage052[246], stage052[247], stage052[248]},
      {stage054[245], stage053[232], stage052[263], stage051[239], stage050[276]}
   );
   gpc615_5 gpc615_5_7637(
      {stage050[263], stage050[264], stage050[265], stage050[266], stage050[267]},
      {stage051[223]},
      {stage052[249], stage052[250], stage052[251], stage052[252], stage052[253], stage052[254]},
      {stage054[246], stage053[233], stage052[264], stage051[240], stage050[277]}
   );
   gpc1_1 gpc1_1_7638(
      {stage051[224]},
      {stage051[241]}
   );
   gpc1_1 gpc1_1_7639(
      {stage051[225]},
      {stage051[242]}
   );
   gpc1_1 gpc1_1_7640(
      {stage051[226]},
      {stage051[243]}
   );
   gpc1_1 gpc1_1_7641(
      {stage051[227]},
      {stage051[244]}
   );
   gpc1_1 gpc1_1_7642(
      {stage051[228]},
      {stage051[245]}
   );
   gpc1_1 gpc1_1_7643(
      {stage051[229]},
      {stage051[246]}
   );
   gpc1_1 gpc1_1_7644(
      {stage051[230]},
      {stage051[247]}
   );
   gpc606_5 gpc606_5_7645(
      {stage051[231], stage051[232], stage051[233], stage051[234], stage051[235], stage051[236]},
      {stage053[212], stage053[213], stage053[214], stage053[215], stage053[216], stage053[217]},
      {stage055[265], stage054[247], stage053[234], stage052[265], stage051[248]}
   );
   gpc1_1 gpc1_1_7646(
      {stage052[255]},
      {stage052[266]}
   );
   gpc1_1 gpc1_1_7647(
      {stage052[256]},
      {stage052[267]}
   );
   gpc1_1 gpc1_1_7648(
      {stage052[257]},
      {stage052[268]}
   );
   gpc1_1 gpc1_1_7649(
      {stage052[258]},
      {stage052[269]}
   );
   gpc1_1 gpc1_1_7650(
      {stage052[259]},
      {stage052[270]}
   );
   gpc1_1 gpc1_1_7651(
      {stage052[260]},
      {stage052[271]}
   );
   gpc1_1 gpc1_1_7652(
      {stage052[261]},
      {stage052[272]}
   );
   gpc1_1 gpc1_1_7653(
      {stage052[262]},
      {stage052[273]}
   );
   gpc1_1 gpc1_1_7654(
      {stage053[218]},
      {stage053[235]}
   );
   gpc1_1 gpc1_1_7655(
      {stage053[219]},
      {stage053[236]}
   );
   gpc1_1 gpc1_1_7656(
      {stage053[220]},
      {stage053[237]}
   );
   gpc1_1 gpc1_1_7657(
      {stage053[221]},
      {stage053[238]}
   );
   gpc1_1 gpc1_1_7658(
      {stage053[222]},
      {stage053[239]}
   );
   gpc1_1 gpc1_1_7659(
      {stage053[223]},
      {stage053[240]}
   );
   gpc1_1 gpc1_1_7660(
      {stage053[224]},
      {stage053[241]}
   );
   gpc1_1 gpc1_1_7661(
      {stage053[225]},
      {stage053[242]}
   );
   gpc1_1 gpc1_1_7662(
      {stage053[226]},
      {stage053[243]}
   );
   gpc1_1 gpc1_1_7663(
      {stage053[227]},
      {stage053[244]}
   );
   gpc1_1 gpc1_1_7664(
      {stage053[228]},
      {stage053[245]}
   );
   gpc1_1 gpc1_1_7665(
      {stage053[229]},
      {stage053[246]}
   );
   gpc1_1 gpc1_1_7666(
      {stage053[230]},
      {stage053[247]}
   );
   gpc1_1 gpc1_1_7667(
      {stage053[231]},
      {stage053[248]}
   );
   gpc1_1 gpc1_1_7668(
      {stage054[234]},
      {stage054[248]}
   );
   gpc1_1 gpc1_1_7669(
      {stage054[235]},
      {stage054[249]}
   );
   gpc1_1 gpc1_1_7670(
      {stage054[236]},
      {stage054[250]}
   );
   gpc1_1 gpc1_1_7671(
      {stage054[237]},
      {stage054[251]}
   );
   gpc1_1 gpc1_1_7672(
      {stage054[238]},
      {stage054[252]}
   );
   gpc1_1 gpc1_1_7673(
      {stage054[239]},
      {stage054[253]}
   );
   gpc615_5 gpc615_5_7674(
      {stage054[240], stage054[241], stage054[242], stage054[243], stage054[244]},
      {stage055[247]},
      {stage056[235], stage056[236], stage056[237], stage056[238], stage056[239], stage056[240]},
      {stage058[222], stage057[246], stage056[263], stage055[266], stage054[254]}
   );
   gpc1_1 gpc1_1_7675(
      {stage055[248]},
      {stage055[267]}
   );
   gpc1_1 gpc1_1_7676(
      {stage055[249]},
      {stage055[268]}
   );
   gpc1_1 gpc1_1_7677(
      {stage055[250]},
      {stage055[269]}
   );
   gpc1_1 gpc1_1_7678(
      {stage055[251]},
      {stage055[270]}
   );
   gpc1_1 gpc1_1_7679(
      {stage055[252]},
      {stage055[271]}
   );
   gpc1_1 gpc1_1_7680(
      {stage055[253]},
      {stage055[272]}
   );
   gpc1_1 gpc1_1_7681(
      {stage055[254]},
      {stage055[273]}
   );
   gpc1_1 gpc1_1_7682(
      {stage055[255]},
      {stage055[274]}
   );
   gpc1_1 gpc1_1_7683(
      {stage055[256]},
      {stage055[275]}
   );
   gpc1_1 gpc1_1_7684(
      {stage055[257]},
      {stage055[276]}
   );
   gpc1_1 gpc1_1_7685(
      {stage055[258]},
      {stage055[277]}
   );
   gpc1_1 gpc1_1_7686(
      {stage055[259]},
      {stage055[278]}
   );
   gpc1_1 gpc1_1_7687(
      {stage055[260]},
      {stage055[279]}
   );
   gpc1_1 gpc1_1_7688(
      {stage055[261]},
      {stage055[280]}
   );
   gpc1_1 gpc1_1_7689(
      {stage055[262]},
      {stage055[281]}
   );
   gpc1_1 gpc1_1_7690(
      {stage055[263]},
      {stage055[282]}
   );
   gpc1_1 gpc1_1_7691(
      {stage055[264]},
      {stage055[283]}
   );
   gpc1_1 gpc1_1_7692(
      {stage056[241]},
      {stage056[264]}
   );
   gpc1_1 gpc1_1_7693(
      {stage056[242]},
      {stage056[265]}
   );
   gpc1_1 gpc1_1_7694(
      {stage056[243]},
      {stage056[266]}
   );
   gpc1_1 gpc1_1_7695(
      {stage056[244]},
      {stage056[267]}
   );
   gpc1_1 gpc1_1_7696(
      {stage056[245]},
      {stage056[268]}
   );
   gpc1_1 gpc1_1_7697(
      {stage056[246]},
      {stage056[269]}
   );
   gpc1_1 gpc1_1_7698(
      {stage056[247]},
      {stage056[270]}
   );
   gpc1_1 gpc1_1_7699(
      {stage056[248]},
      {stage056[271]}
   );
   gpc1_1 gpc1_1_7700(
      {stage056[249]},
      {stage056[272]}
   );
   gpc1_1 gpc1_1_7701(
      {stage056[250]},
      {stage056[273]}
   );
   gpc1_1 gpc1_1_7702(
      {stage056[251]},
      {stage056[274]}
   );
   gpc1_1 gpc1_1_7703(
      {stage056[252]},
      {stage056[275]}
   );
   gpc1_1 gpc1_1_7704(
      {stage056[253]},
      {stage056[276]}
   );
   gpc1_1 gpc1_1_7705(
      {stage056[254]},
      {stage056[277]}
   );
   gpc1_1 gpc1_1_7706(
      {stage056[255]},
      {stage056[278]}
   );
   gpc1_1 gpc1_1_7707(
      {stage056[256]},
      {stage056[279]}
   );
   gpc1_1 gpc1_1_7708(
      {stage056[257]},
      {stage056[280]}
   );
   gpc1_1 gpc1_1_7709(
      {stage056[258]},
      {stage056[281]}
   );
   gpc1_1 gpc1_1_7710(
      {stage056[259]},
      {stage056[282]}
   );
   gpc1_1 gpc1_1_7711(
      {stage056[260]},
      {stage056[283]}
   );
   gpc1_1 gpc1_1_7712(
      {stage056[261]},
      {stage056[284]}
   );
   gpc1_1 gpc1_1_7713(
      {stage056[262]},
      {stage056[285]}
   );
   gpc1_1 gpc1_1_7714(
      {stage057[233]},
      {stage057[247]}
   );
   gpc1_1 gpc1_1_7715(
      {stage057[234]},
      {stage057[248]}
   );
   gpc1_1 gpc1_1_7716(
      {stage057[235]},
      {stage057[249]}
   );
   gpc615_5 gpc615_5_7717(
      {stage057[236], stage057[237], stage057[238], stage057[239], stage057[240]},
      {stage058[209]},
      {stage059[267], stage059[268], stage059[269], stage059[270], stage059[271], stage059[272]},
      {stage061[262], stage060[229], stage059[297], stage058[223], stage057[250]}
   );
   gpc615_5 gpc615_5_7718(
      {stage057[241], stage057[242], stage057[243], stage057[244], stage057[245]},
      {stage058[210]},
      {stage059[273], stage059[274], stage059[275], stage059[276], stage059[277], stage059[278]},
      {stage061[263], stage060[230], stage059[298], stage058[224], stage057[251]}
   );
   gpc1_1 gpc1_1_7719(
      {stage058[211]},
      {stage058[225]}
   );
   gpc1_1 gpc1_1_7720(
      {stage058[212]},
      {stage058[226]}
   );
   gpc1_1 gpc1_1_7721(
      {stage058[213]},
      {stage058[227]}
   );
   gpc1_1 gpc1_1_7722(
      {stage058[214]},
      {stage058[228]}
   );
   gpc1_1 gpc1_1_7723(
      {stage058[215]},
      {stage058[229]}
   );
   gpc1_1 gpc1_1_7724(
      {stage058[216]},
      {stage058[230]}
   );
   gpc615_5 gpc615_5_7725(
      {stage058[217], stage058[218], stage058[219], stage058[220], stage058[221]},
      {stage059[279]},
      {stage060[215], stage060[216], stage060[217], stage060[218], stage060[219], stage060[220]},
      {stage062[239], stage061[264], stage060[231], stage059[299], stage058[231]}
   );
   gpc1_1 gpc1_1_7726(
      {stage059[280]},
      {stage059[300]}
   );
   gpc1_1 gpc1_1_7727(
      {stage059[281]},
      {stage059[301]}
   );
   gpc1_1 gpc1_1_7728(
      {stage059[282]},
      {stage059[302]}
   );
   gpc1_1 gpc1_1_7729(
      {stage059[283]},
      {stage059[303]}
   );
   gpc1_1 gpc1_1_7730(
      {stage059[284]},
      {stage059[304]}
   );
   gpc1_1 gpc1_1_7731(
      {stage059[285]},
      {stage059[305]}
   );
   gpc1_1 gpc1_1_7732(
      {stage059[286]},
      {stage059[306]}
   );
   gpc1_1 gpc1_1_7733(
      {stage059[287]},
      {stage059[307]}
   );
   gpc1_1 gpc1_1_7734(
      {stage059[288]},
      {stage059[308]}
   );
   gpc1_1 gpc1_1_7735(
      {stage059[289]},
      {stage059[309]}
   );
   gpc1_1 gpc1_1_7736(
      {stage059[290]},
      {stage059[310]}
   );
   gpc1_1 gpc1_1_7737(
      {stage059[291]},
      {stage059[311]}
   );
   gpc615_5 gpc615_5_7738(
      {stage059[292], stage059[293], stage059[294], stage059[295], stage059[296]},
      {stage060[221]},
      {stage061[246], stage061[247], stage061[248], stage061[249], stage061[250], stage061[251]},
      {stage063[209], stage062[240], stage061[265], stage060[232], stage059[312]}
   );
   gpc1_1 gpc1_1_7739(
      {stage060[222]},
      {stage060[233]}
   );
   gpc1_1 gpc1_1_7740(
      {stage060[223]},
      {stage060[234]}
   );
   gpc1_1 gpc1_1_7741(
      {stage060[224]},
      {stage060[235]}
   );
   gpc1_1 gpc1_1_7742(
      {stage060[225]},
      {stage060[236]}
   );
   gpc1_1 gpc1_1_7743(
      {stage060[226]},
      {stage060[237]}
   );
   gpc1_1 gpc1_1_7744(
      {stage060[227]},
      {stage060[238]}
   );
   gpc1_1 gpc1_1_7745(
      {stage060[228]},
      {stage060[239]}
   );
   gpc1_1 gpc1_1_7746(
      {stage061[252]},
      {stage061[266]}
   );
   gpc1_1 gpc1_1_7747(
      {stage061[253]},
      {stage061[267]}
   );
   gpc1_1 gpc1_1_7748(
      {stage061[254]},
      {stage061[268]}
   );
   gpc1_1 gpc1_1_7749(
      {stage061[255]},
      {stage061[269]}
   );
   gpc1_1 gpc1_1_7750(
      {stage061[256]},
      {stage061[270]}
   );
   gpc1_1 gpc1_1_7751(
      {stage061[257]},
      {stage061[271]}
   );
   gpc1_1 gpc1_1_7752(
      {stage061[258]},
      {stage061[272]}
   );
   gpc1_1 gpc1_1_7753(
      {stage061[259]},
      {stage061[273]}
   );
   gpc1_1 gpc1_1_7754(
      {stage061[260]},
      {stage061[274]}
   );
   gpc1_1 gpc1_1_7755(
      {stage061[261]},
      {stage061[275]}
   );
   gpc1_1 gpc1_1_7756(
      {stage062[215]},
      {stage062[241]}
   );
   gpc1_1 gpc1_1_7757(
      {stage062[216]},
      {stage062[242]}
   );
   gpc1_1 gpc1_1_7758(
      {stage062[217]},
      {stage062[243]}
   );
   gpc1_1 gpc1_1_7759(
      {stage062[218]},
      {stage062[244]}
   );
   gpc1_1 gpc1_1_7760(
      {stage062[219]},
      {stage062[245]}
   );
   gpc1_1 gpc1_1_7761(
      {stage062[220]},
      {stage062[246]}
   );
   gpc1_1 gpc1_1_7762(
      {stage062[221]},
      {stage062[247]}
   );
   gpc1_1 gpc1_1_7763(
      {stage062[222]},
      {stage062[248]}
   );
   gpc1_1 gpc1_1_7764(
      {stage062[223]},
      {stage062[249]}
   );
   gpc1_1 gpc1_1_7765(
      {stage062[224]},
      {stage062[250]}
   );
   gpc207_4 gpc207_4_7766(
      {stage062[225], stage062[226], stage062[227], stage062[228], stage062[229], stage062[230], stage062[231]},
      {stage064[244], stage064[245]},
      {stage065[255], stage064[257], stage063[210], stage062[251]}
   );
   gpc207_4 gpc207_4_7767(
      {stage062[232], stage062[233], stage062[234], stage062[235], stage062[236], stage062[237], stage062[238]},
      {stage064[246], stage064[247]},
      {stage065[256], stage064[258], stage063[211], stage062[252]}
   );
   gpc606_5 gpc606_5_7768(
      {stage063[193], stage063[194], stage063[195], stage063[196], stage063[197], stage063[198]},
      {stage065[237], stage065[238], stage065[239], stage065[240], stage065[241], stage065[242]},
      {stage067[253], stage066[273], stage065[257], stage064[259], stage063[212]}
   );
   gpc615_5 gpc615_5_7769(
      {stage063[199], stage063[200], stage063[201], stage063[202], stage063[203]},
      {stage064[248]},
      {stage065[243], stage065[244], stage065[245], stage065[246], stage065[247], stage065[248]},
      {stage067[254], stage066[274], stage065[258], stage064[260], stage063[213]}
   );
   gpc615_5 gpc615_5_7770(
      {stage063[204], stage063[205], stage063[206], stage063[207], stage063[208]},
      {stage064[249]},
      {stage065[249], stage065[250], stage065[251], stage065[252], stage065[253], stage065[254]},
      {stage067[255], stage066[275], stage065[259], stage064[261], stage063[214]}
   );
   gpc1_1 gpc1_1_7771(
      {stage064[250]},
      {stage064[262]}
   );
   gpc606_5 gpc606_5_7772(
      {stage064[251], stage064[252], stage064[253], stage064[254], stage064[255], stage064[256]},
      {stage066[246], stage066[247], stage066[248], stage066[249], stage066[250], stage066[251]},
      {stage068[266], stage067[256], stage066[276], stage065[260], stage064[263]}
   );
   gpc1_1 gpc1_1_7773(
      {stage066[252]},
      {stage066[277]}
   );
   gpc1_1 gpc1_1_7774(
      {stage066[253]},
      {stage066[278]}
   );
   gpc1_1 gpc1_1_7775(
      {stage066[254]},
      {stage066[279]}
   );
   gpc1_1 gpc1_1_7776(
      {stage066[255]},
      {stage066[280]}
   );
   gpc1_1 gpc1_1_7777(
      {stage066[256]},
      {stage066[281]}
   );
   gpc1_1 gpc1_1_7778(
      {stage066[257]},
      {stage066[282]}
   );
   gpc615_5 gpc615_5_7779(
      {stage066[258], stage066[259], stage066[260], stage066[261], stage066[262]},
      {stage067[244]},
      {stage068[241], stage068[242], stage068[243], stage068[244], stage068[245], stage068[246]},
      {stage070[249], stage069[256], stage068[267], stage067[257], stage066[283]}
   );
   gpc615_5 gpc615_5_7780(
      {stage066[263], stage066[264], stage066[265], stage066[266], stage066[267]},
      {stage067[245]},
      {stage068[247], stage068[248], stage068[249], stage068[250], stage068[251], stage068[252]},
      {stage070[250], stage069[257], stage068[268], stage067[258], stage066[284]}
   );
   gpc615_5 gpc615_5_7781(
      {stage066[268], stage066[269], stage066[270], stage066[271], stage066[272]},
      {stage067[246]},
      {stage068[253], stage068[254], stage068[255], stage068[256], stage068[257], stage068[258]},
      {stage070[251], stage069[258], stage068[269], stage067[259], stage066[285]}
   );
   gpc1_1 gpc1_1_7782(
      {stage067[247]},
      {stage067[260]}
   );
   gpc615_5 gpc615_5_7783(
      {stage067[248], stage067[249], stage067[250], stage067[251], stage067[252]},
      {stage068[259]},
      {stage069[233], stage069[234], stage069[235], stage069[236], stage069[237], stage069[238]},
      {stage071[256], stage070[252], stage069[259], stage068[270], stage067[261]}
   );
   gpc1_1 gpc1_1_7784(
      {stage068[260]},
      {stage068[271]}
   );
   gpc1_1 gpc1_1_7785(
      {stage068[261]},
      {stage068[272]}
   );
   gpc1_1 gpc1_1_7786(
      {stage068[262]},
      {stage068[273]}
   );
   gpc1_1 gpc1_1_7787(
      {stage068[263]},
      {stage068[274]}
   );
   gpc1_1 gpc1_1_7788(
      {stage068[264]},
      {stage068[275]}
   );
   gpc1_1 gpc1_1_7789(
      {stage068[265]},
      {stage068[276]}
   );
   gpc606_5 gpc606_5_7790(
      {stage069[239], stage069[240], stage069[241], stage069[242], stage069[243], stage069[244]},
      {stage071[237], stage071[238], stage071[239], stage071[240], stage071[241], stage071[242]},
      {stage073[232], stage072[299], stage071[257], stage070[253], stage069[260]}
   );
   gpc606_5 gpc606_5_7791(
      {stage069[245], stage069[246], stage069[247], stage069[248], stage069[249], stage069[250]},
      {stage071[243], stage071[244], stage071[245], stage071[246], stage071[247], stage071[248]},
      {stage073[233], stage072[300], stage071[258], stage070[254], stage069[261]}
   );
   gpc606_5 gpc606_5_7792(
      {stage069[251], stage069[252], stage069[253], stage069[254], stage069[255], 1'h0},
      {stage071[249], stage071[250], stage071[251], stage071[252], stage071[253], stage071[254]},
      {stage073[234], stage072[301], stage071[259], stage070[255], stage069[262]}
   );
   gpc615_5 gpc615_5_7793(
      {stage070[234], stage070[235], stage070[236], stage070[237], stage070[238]},
      {stage071[255]},
      {stage072[267], stage072[268], stage072[269], stage072[270], stage072[271], stage072[272]},
      {stage074[243], stage073[235], stage072[302], stage071[260], stage070[256]}
   );
   gpc615_5 gpc615_5_7794(
      {stage070[239], stage070[240], stage070[241], stage070[242], stage070[243]},
      {1'h0},
      {stage072[273], stage072[274], stage072[275], stage072[276], stage072[277], stage072[278]},
      {stage074[244], stage073[236], stage072[303], stage071[261], stage070[257]}
   );
   gpc615_5 gpc615_5_7795(
      {stage070[244], stage070[245], stage070[246], stage070[247], stage070[248]},
      {1'h0},
      {stage072[279], stage072[280], stage072[281], stage072[282], stage072[283], stage072[284]},
      {stage074[245], stage073[237], stage072[304], stage071[262], stage070[258]}
   );
   gpc1_1 gpc1_1_7796(
      {stage072[285]},
      {stage072[305]}
   );
   gpc1_1 gpc1_1_7797(
      {stage072[286]},
      {stage072[306]}
   );
   gpc1_1 gpc1_1_7798(
      {stage072[287]},
      {stage072[307]}
   );
   gpc1_1 gpc1_1_7799(
      {stage072[288]},
      {stage072[308]}
   );
   gpc615_5 gpc615_5_7800(
      {stage072[289], stage072[290], stage072[291], stage072[292], stage072[293]},
      {stage073[217]},
      {stage074[227], stage074[228], stage074[229], stage074[230], stage074[231], stage074[232]},
      {stage076[209], stage075[205], stage074[246], stage073[238], stage072[309]}
   );
   gpc615_5 gpc615_5_7801(
      {stage072[294], stage072[295], stage072[296], stage072[297], stage072[298]},
      {stage073[218]},
      {stage074[233], stage074[234], stage074[235], stage074[236], stage074[237], stage074[238]},
      {stage076[210], stage075[206], stage074[247], stage073[239], stage072[310]}
   );
   gpc1_1 gpc1_1_7802(
      {stage073[219]},
      {stage073[240]}
   );
   gpc606_5 gpc606_5_7803(
      {stage073[220], stage073[221], stage073[222], stage073[223], stage073[224], stage073[225]},
      {stage075[193], stage075[194], stage075[195], stage075[196], stage075[197], stage075[198]},
      {stage077[243], stage076[211], stage075[207], stage074[248], stage073[241]}
   );
   gpc606_5 gpc606_5_7804(
      {stage073[226], stage073[227], stage073[228], stage073[229], stage073[230], stage073[231]},
      {stage075[199], stage075[200], stage075[201], stage075[202], stage075[203], stage075[204]},
      {stage077[244], stage076[212], stage075[208], stage074[249], stage073[242]}
   );
   gpc1_1 gpc1_1_7805(
      {stage074[239]},
      {stage074[250]}
   );
   gpc1_1 gpc1_1_7806(
      {stage074[240]},
      {stage074[251]}
   );
   gpc1_1 gpc1_1_7807(
      {stage074[241]},
      {stage074[252]}
   );
   gpc1_1 gpc1_1_7808(
      {stage074[242]},
      {stage074[253]}
   );
   gpc615_5 gpc615_5_7809(
      {stage076[197], stage076[198], stage076[199], stage076[200], stage076[201]},
      {stage077[230]},
      {stage078[207], stage078[208], stage078[209], stage078[210], stage078[211], stage078[212]},
      {stage080[253], stage079[238], stage078[228], stage077[245], stage076[213]}
   );
   gpc207_4 gpc207_4_7810(
      {stage076[202], stage076[203], stage076[204], stage076[205], stage076[206], stage076[207], stage076[208]},
      {stage078[213], stage078[214]},
      {stage079[239], stage078[229], stage077[246], stage076[214]}
   );
   gpc1_1 gpc1_1_7811(
      {stage077[231]},
      {stage077[247]}
   );
   gpc1_1 gpc1_1_7812(
      {stage077[232]},
      {stage077[248]}
   );
   gpc1_1 gpc1_1_7813(
      {stage077[233]},
      {stage077[249]}
   );
   gpc623_5 gpc623_5_7814(
      {stage077[234], stage077[235], stage077[236]},
      {stage078[215], stage078[216]},
      {stage079[216], stage079[217], stage079[218], stage079[219], stage079[220], stage079[221]},
      {stage081[258], stage080[254], stage079[240], stage078[230], stage077[250]}
   );
   gpc606_5 gpc606_5_7815(
      {stage077[237], stage077[238], stage077[239], stage077[240], stage077[241], stage077[242]},
      {stage079[222], stage079[223], stage079[224], stage079[225], stage079[226], stage079[227]},
      {stage081[259], stage080[255], stage079[241], stage078[231], stage077[251]}
   );
   gpc606_5 gpc606_5_7816(
      {stage078[217], stage078[218], stage078[219], stage078[220], stage078[221], stage078[222]},
      {stage080[232], stage080[233], stage080[234], stage080[235], stage080[236], stage080[237]},
      {stage082[255], stage081[260], stage080[256], stage079[242], stage078[232]}
   );
   gpc615_5 gpc615_5_7817(
      {stage078[223], stage078[224], stage078[225], stage078[226], stage078[227]},
      {stage079[228]},
      {stage080[238], stage080[239], stage080[240], stage080[241], stage080[242], stage080[243]},
      {stage082[256], stage081[261], stage080[257], stage079[243], stage078[233]}
   );
   gpc1_1 gpc1_1_7818(
      {stage079[229]},
      {stage079[244]}
   );
   gpc1_1 gpc1_1_7819(
      {stage079[230]},
      {stage079[245]}
   );
   gpc1_1 gpc1_1_7820(
      {stage079[231]},
      {stage079[246]}
   );
   gpc1_1 gpc1_1_7821(
      {stage079[232]},
      {stage079[247]}
   );
   gpc1_1 gpc1_1_7822(
      {stage079[233]},
      {stage079[248]}
   );
   gpc1_1 gpc1_1_7823(
      {stage079[234]},
      {stage079[249]}
   );
   gpc1_1 gpc1_1_7824(
      {stage079[235]},
      {stage079[250]}
   );
   gpc1_1 gpc1_1_7825(
      {stage079[236]},
      {stage079[251]}
   );
   gpc1_1 gpc1_1_7826(
      {stage079[237]},
      {stage079[252]}
   );
   gpc1_1 gpc1_1_7827(
      {stage080[244]},
      {stage080[258]}
   );
   gpc1_1 gpc1_1_7828(
      {stage080[245]},
      {stage080[259]}
   );
   gpc7_3 gpc7_3_7829(
      {stage080[246], stage080[247], stage080[248], stage080[249], stage080[250], stage080[251], stage080[252]},
      {stage082[257], stage081[262], stage080[260]}
   );
   gpc1_1 gpc1_1_7830(
      {stage081[238]},
      {stage081[263]}
   );
   gpc1_1 gpc1_1_7831(
      {stage081[239]},
      {stage081[264]}
   );
   gpc1_1 gpc1_1_7832(
      {stage081[240]},
      {stage081[265]}
   );
   gpc1_1 gpc1_1_7833(
      {stage081[241]},
      {stage081[266]}
   );
   gpc1_1 gpc1_1_7834(
      {stage081[242]},
      {stage081[267]}
   );
   gpc1_1 gpc1_1_7835(
      {stage081[243]},
      {stage081[268]}
   );
   gpc1_1 gpc1_1_7836(
      {stage081[244]},
      {stage081[269]}
   );
   gpc1_1 gpc1_1_7837(
      {stage081[245]},
      {stage081[270]}
   );
   gpc1_1 gpc1_1_7838(
      {stage081[246]},
      {stage081[271]}
   );
   gpc1_1 gpc1_1_7839(
      {stage081[247]},
      {stage081[272]}
   );
   gpc1_1 gpc1_1_7840(
      {stage081[248]},
      {stage081[273]}
   );
   gpc1_1 gpc1_1_7841(
      {stage081[249]},
      {stage081[274]}
   );
   gpc1_1 gpc1_1_7842(
      {stage081[250]},
      {stage081[275]}
   );
   gpc1_1 gpc1_1_7843(
      {stage081[251]},
      {stage081[276]}
   );
   gpc1_1 gpc1_1_7844(
      {stage081[252]},
      {stage081[277]}
   );
   gpc1_1 gpc1_1_7845(
      {stage081[253]},
      {stage081[278]}
   );
   gpc1_1 gpc1_1_7846(
      {stage081[254]},
      {stage081[279]}
   );
   gpc1_1 gpc1_1_7847(
      {stage081[255]},
      {stage081[280]}
   );
   gpc1_1 gpc1_1_7848(
      {stage081[256]},
      {stage081[281]}
   );
   gpc1_1 gpc1_1_7849(
      {stage081[257]},
      {stage081[282]}
   );
   gpc1_1 gpc1_1_7850(
      {stage082[240]},
      {stage082[258]}
   );
   gpc1_1 gpc1_1_7851(
      {stage082[241]},
      {stage082[259]}
   );
   gpc1_1 gpc1_1_7852(
      {stage082[242]},
      {stage082[260]}
   );
   gpc606_5 gpc606_5_7853(
      {stage082[243], stage082[244], stage082[245], stage082[246], stage082[247], stage082[248]},
      {stage084[218], stage084[219], stage084[220], stage084[221], stage084[222], stage084[223]},
      {stage086[271], stage085[265], stage084[235], stage083[261], stage082[261]}
   );
   gpc606_5 gpc606_5_7854(
      {stage082[249], stage082[250], stage082[251], stage082[252], stage082[253], stage082[254]},
      {stage084[224], stage084[225], stage084[226], stage084[227], stage084[228], stage084[229]},
      {stage086[272], stage085[266], stage084[236], stage083[262], stage082[262]}
   );
   gpc1_1 gpc1_1_7855(
      {stage083[246]},
      {stage083[263]}
   );
   gpc1_1 gpc1_1_7856(
      {stage083[247]},
      {stage083[264]}
   );
   gpc1_1 gpc1_1_7857(
      {stage083[248]},
      {stage083[265]}
   );
   gpc606_5 gpc606_5_7858(
      {stage083[249], stage083[250], stage083[251], stage083[252], stage083[253], stage083[254]},
      {stage085[249], stage085[250], stage085[251], stage085[252], stage085[253], stage085[254]},
      {stage087[223], stage086[273], stage085[267], stage084[237], stage083[266]}
   );
   gpc606_5 gpc606_5_7859(
      {stage083[255], stage083[256], stage083[257], stage083[258], stage083[259], stage083[260]},
      {stage085[255], stage085[256], stage085[257], stage085[258], stage085[259], stage085[260]},
      {stage087[224], stage086[274], stage085[268], stage084[238], stage083[267]}
   );
   gpc606_5 gpc606_5_7860(
      {stage084[230], stage084[231], stage084[232], stage084[233], stage084[234], 1'h0},
      {stage086[243], stage086[244], stage086[245], stage086[246], stage086[247], stage086[248]},
      {stage088[264], stage087[225], stage086[275], stage085[269], stage084[239]}
   );
   gpc1_1 gpc1_1_7861(
      {stage085[261]},
      {stage085[270]}
   );
   gpc1_1 gpc1_1_7862(
      {stage085[262]},
      {stage085[271]}
   );
   gpc1_1 gpc1_1_7863(
      {stage085[263]},
      {stage085[272]}
   );
   gpc1_1 gpc1_1_7864(
      {stage085[264]},
      {stage085[273]}
   );
   gpc1_1 gpc1_1_7865(
      {stage086[249]},
      {stage086[276]}
   );
   gpc1_1 gpc1_1_7866(
      {stage086[250]},
      {stage086[277]}
   );
   gpc1_1 gpc1_1_7867(
      {stage086[251]},
      {stage086[278]}
   );
   gpc1_1 gpc1_1_7868(
      {stage086[252]},
      {stage086[279]}
   );
   gpc1_1 gpc1_1_7869(
      {stage086[253]},
      {stage086[280]}
   );
   gpc7_3 gpc7_3_7870(
      {stage086[254], stage086[255], stage086[256], stage086[257], stage086[258], stage086[259], stage086[260]},
      {stage088[265], stage087[226], stage086[281]}
   );
   gpc615_5 gpc615_5_7871(
      {stage086[261], stage086[262], stage086[263], stage086[264], stage086[265]},
      {stage087[213]},
      {stage088[246], stage088[247], stage088[248], stage088[249], stage088[250], stage088[251]},
      {stage090[231], stage089[247], stage088[266], stage087[227], stage086[282]}
   );
   gpc615_5 gpc615_5_7872(
      {stage086[266], stage086[267], stage086[268], stage086[269], stage086[270]},
      {stage087[214]},
      {stage088[252], stage088[253], stage088[254], stage088[255], stage088[256], stage088[257]},
      {stage090[232], stage089[248], stage088[267], stage087[228], stage086[283]}
   );
   gpc1_1 gpc1_1_7873(
      {stage087[215]},
      {stage087[229]}
   );
   gpc1_1 gpc1_1_7874(
      {stage087[216]},
      {stage087[230]}
   );
   gpc1_1 gpc1_1_7875(
      {stage087[217]},
      {stage087[231]}
   );
   gpc1_1 gpc1_1_7876(
      {stage087[218]},
      {stage087[232]}
   );
   gpc1_1 gpc1_1_7877(
      {stage087[219]},
      {stage087[233]}
   );
   gpc1_1 gpc1_1_7878(
      {stage087[220]},
      {stage087[234]}
   );
   gpc1_1 gpc1_1_7879(
      {stage087[221]},
      {stage087[235]}
   );
   gpc1_1 gpc1_1_7880(
      {stage087[222]},
      {stage087[236]}
   );
   gpc1_1 gpc1_1_7881(
      {stage088[258]},
      {stage088[268]}
   );
   gpc1_1 gpc1_1_7882(
      {stage088[259]},
      {stage088[269]}
   );
   gpc1_1 gpc1_1_7883(
      {stage088[260]},
      {stage088[270]}
   );
   gpc1_1 gpc1_1_7884(
      {stage088[261]},
      {stage088[271]}
   );
   gpc1_1 gpc1_1_7885(
      {stage088[262]},
      {stage088[272]}
   );
   gpc1_1 gpc1_1_7886(
      {stage088[263]},
      {stage088[273]}
   );
   gpc1_1 gpc1_1_7887(
      {stage089[216]},
      {stage089[249]}
   );
   gpc1_1 gpc1_1_7888(
      {stage089[217]},
      {stage089[250]}
   );
   gpc1_1 gpc1_1_7889(
      {stage089[218]},
      {stage089[251]}
   );
   gpc1_1 gpc1_1_7890(
      {stage089[219]},
      {stage089[252]}
   );
   gpc1_1 gpc1_1_7891(
      {stage089[220]},
      {stage089[253]}
   );
   gpc1_1 gpc1_1_7892(
      {stage089[221]},
      {stage089[254]}
   );
   gpc1_1 gpc1_1_7893(
      {stage089[222]},
      {stage089[255]}
   );
   gpc1_1 gpc1_1_7894(
      {stage089[223]},
      {stage089[256]}
   );
   gpc1_1 gpc1_1_7895(
      {stage089[224]},
      {stage089[257]}
   );
   gpc1_1 gpc1_1_7896(
      {stage089[225]},
      {stage089[258]}
   );
   gpc1_1 gpc1_1_7897(
      {stage089[226]},
      {stage089[259]}
   );
   gpc1_1 gpc1_1_7898(
      {stage089[227]},
      {stage089[260]}
   );
   gpc1_1 gpc1_1_7899(
      {stage089[228]},
      {stage089[261]}
   );
   gpc1_1 gpc1_1_7900(
      {stage089[229]},
      {stage089[262]}
   );
   gpc606_5 gpc606_5_7901(
      {stage089[230], stage089[231], stage089[232], stage089[233], stage089[234], stage089[235]},
      {stage091[255], stage091[256], stage091[257], stage091[258], stage091[259], stage091[260]},
      {stage093[221], stage092[241], stage091[302], stage090[233], stage089[263]}
   );
   gpc606_5 gpc606_5_7902(
      {stage089[236], stage089[237], stage089[238], stage089[239], stage089[240], stage089[241]},
      {stage091[261], stage091[262], stage091[263], stage091[264], stage091[265], stage091[266]},
      {stage093[222], stage092[242], stage091[303], stage090[234], stage089[264]}
   );
   gpc615_5 gpc615_5_7903(
      {stage089[242], stage089[243], stage089[244], stage089[245], stage089[246]},
      {stage090[217]},
      {stage091[267], stage091[268], stage091[269], stage091[270], stage091[271], stage091[272]},
      {stage093[223], stage092[243], stage091[304], stage090[235], stage089[265]}
   );
   gpc1_1 gpc1_1_7904(
      {stage090[218]},
      {stage090[236]}
   );
   gpc1_1 gpc1_1_7905(
      {stage090[219]},
      {stage090[237]}
   );
   gpc1_1 gpc1_1_7906(
      {stage090[220]},
      {stage090[238]}
   );
   gpc1_1 gpc1_1_7907(
      {stage090[221]},
      {stage090[239]}
   );
   gpc1_1 gpc1_1_7908(
      {stage090[222]},
      {stage090[240]}
   );
   gpc1_1 gpc1_1_7909(
      {stage090[223]},
      {stage090[241]}
   );
   gpc1_1 gpc1_1_7910(
      {stage090[224]},
      {stage090[242]}
   );
   gpc1_1 gpc1_1_7911(
      {stage090[225]},
      {stage090[243]}
   );
   gpc615_5 gpc615_5_7912(
      {stage090[226], stage090[227], stage090[228], stage090[229], stage090[230]},
      {stage091[273]},
      {stage092[227], stage092[228], stage092[229], stage092[230], stage092[231], stage092[232]},
      {stage094[236], stage093[224], stage092[244], stage091[305], stage090[244]}
   );
   gpc1_1 gpc1_1_7913(
      {stage091[274]},
      {stage091[306]}
   );
   gpc1_1 gpc1_1_7914(
      {stage091[275]},
      {stage091[307]}
   );
   gpc1_1 gpc1_1_7915(
      {stage091[276]},
      {stage091[308]}
   );
   gpc1_1 gpc1_1_7916(
      {stage091[277]},
      {stage091[309]}
   );
   gpc1_1 gpc1_1_7917(
      {stage091[278]},
      {stage091[310]}
   );
   gpc1_1 gpc1_1_7918(
      {stage091[279]},
      {stage091[311]}
   );
   gpc1_1 gpc1_1_7919(
      {stage091[280]},
      {stage091[312]}
   );
   gpc1_1 gpc1_1_7920(
      {stage091[281]},
      {stage091[313]}
   );
   gpc1_1 gpc1_1_7921(
      {stage091[282]},
      {stage091[314]}
   );
   gpc1_1 gpc1_1_7922(
      {stage091[283]},
      {stage091[315]}
   );
   gpc1_1 gpc1_1_7923(
      {stage091[284]},
      {stage091[316]}
   );
   gpc1_1 gpc1_1_7924(
      {stage091[285]},
      {stage091[317]}
   );
   gpc1_1 gpc1_1_7925(
      {stage091[286]},
      {stage091[318]}
   );
   gpc1_1 gpc1_1_7926(
      {stage091[287]},
      {stage091[319]}
   );
   gpc1_1 gpc1_1_7927(
      {stage091[288]},
      {stage091[320]}
   );
   gpc1_1 gpc1_1_7928(
      {stage091[289]},
      {stage091[321]}
   );
   gpc1_1 gpc1_1_7929(
      {stage091[290]},
      {stage091[322]}
   );
   gpc1_1 gpc1_1_7930(
      {stage091[291]},
      {stage091[323]}
   );
   gpc1_1 gpc1_1_7931(
      {stage091[292]},
      {stage091[324]}
   );
   gpc1_1 gpc1_1_7932(
      {stage091[293]},
      {stage091[325]}
   );
   gpc1_1 gpc1_1_7933(
      {stage091[294]},
      {stage091[326]}
   );
   gpc1_1 gpc1_1_7934(
      {stage091[295]},
      {stage091[327]}
   );
   gpc1_1 gpc1_1_7935(
      {stage091[296]},
      {stage091[328]}
   );
   gpc615_5 gpc615_5_7936(
      {stage091[297], stage091[298], stage091[299], stage091[300], stage091[301]},
      {stage092[233]},
      {stage093[209], stage093[210], stage093[211], stage093[212], stage093[213], stage093[214]},
      {stage095[214], stage094[237], stage093[225], stage092[245], stage091[329]}
   );
   gpc1_1 gpc1_1_7937(
      {stage092[234]},
      {stage092[246]}
   );
   gpc606_5 gpc606_5_7938(
      {stage092[235], stage092[236], stage092[237], stage092[238], stage092[239], stage092[240]},
      {stage094[224], stage094[225], stage094[226], stage094[227], stage094[228], stage094[229]},
      {stage096[231], stage095[215], stage094[238], stage093[226], stage092[247]}
   );
   gpc1_1 gpc1_1_7939(
      {stage093[215]},
      {stage093[227]}
   );
   gpc1_1 gpc1_1_7940(
      {stage093[216]},
      {stage093[228]}
   );
   gpc1_1 gpc1_1_7941(
      {stage093[217]},
      {stage093[229]}
   );
   gpc1_1 gpc1_1_7942(
      {stage093[218]},
      {stage093[230]}
   );
   gpc1_1 gpc1_1_7943(
      {stage093[219]},
      {stage093[231]}
   );
   gpc1_1 gpc1_1_7944(
      {stage093[220]},
      {stage093[232]}
   );
   gpc606_5 gpc606_5_7945(
      {stage094[230], stage094[231], stage094[232], stage094[233], stage094[234], stage094[235]},
      {stage096[218], stage096[219], stage096[220], stage096[221], stage096[222], stage096[223]},
      {stage098[226], stage097[220], stage096[232], stage095[216], stage094[239]}
   );
   gpc1_1 gpc1_1_7946(
      {stage095[205]},
      {stage095[217]}
   );
   gpc1_1 gpc1_1_7947(
      {stage095[206]},
      {stage095[218]}
   );
   gpc1_1 gpc1_1_7948(
      {stage095[207]},
      {stage095[219]}
   );
   gpc606_5 gpc606_5_7949(
      {stage095[208], stage095[209], stage095[210], stage095[211], stage095[212], stage095[213]},
      {stage097[205], stage097[206], stage097[207], stage097[208], stage097[209], stage097[210]},
      {stage099[280], stage098[227], stage097[221], stage096[233], stage095[220]}
   );
   gpc1_1 gpc1_1_7950(
      {stage096[224]},
      {stage096[234]}
   );
   gpc1_1 gpc1_1_7951(
      {stage096[225]},
      {stage096[235]}
   );
   gpc1_1 gpc1_1_7952(
      {stage096[226]},
      {stage096[236]}
   );
   gpc1_1 gpc1_1_7953(
      {stage096[227]},
      {stage096[237]}
   );
   gpc1_1 gpc1_1_7954(
      {stage096[228]},
      {stage096[238]}
   );
   gpc1_1 gpc1_1_7955(
      {stage096[229]},
      {stage096[239]}
   );
   gpc1_1 gpc1_1_7956(
      {stage096[230]},
      {stage096[240]}
   );
   gpc1_1 gpc1_1_7957(
      {stage097[211]},
      {stage097[222]}
   );
   gpc1_1 gpc1_1_7958(
      {stage097[212]},
      {stage097[223]}
   );
   gpc7_3 gpc7_3_7959(
      {stage097[213], stage097[214], stage097[215], stage097[216], stage097[217], stage097[218], stage097[219]},
      {stage099[281], stage098[228], stage097[224]}
   );
   gpc1_1 gpc1_1_7960(
      {stage098[206]},
      {stage098[229]}
   );
   gpc1_1 gpc1_1_7961(
      {stage098[207]},
      {stage098[230]}
   );
   gpc1_1 gpc1_1_7962(
      {stage098[208]},
      {stage098[231]}
   );
   gpc1_1 gpc1_1_7963(
      {stage098[209]},
      {stage098[232]}
   );
   gpc1_1 gpc1_1_7964(
      {stage098[210]},
      {stage098[233]}
   );
   gpc1_1 gpc1_1_7965(
      {stage098[211]},
      {stage098[234]}
   );
   gpc1_1 gpc1_1_7966(
      {stage098[212]},
      {stage098[235]}
   );
   gpc1_1 gpc1_1_7967(
      {stage098[213]},
      {stage098[236]}
   );
   gpc7_3 gpc7_3_7968(
      {stage098[214], stage098[215], stage098[216], stage098[217], stage098[218], stage098[219], stage098[220]},
      {stage100[218], stage099[282], stage098[237]}
   );
   gpc615_5 gpc615_5_7969(
      {stage098[221], stage098[222], stage098[223], stage098[224], stage098[225]},
      {stage099[258]},
      {stage100[202], stage100[203], stage100[204], stage100[205], stage100[206], stage100[207]},
      {stage102[235], stage101[253], stage100[219], stage099[283], stage098[238]}
   );
   gpc1_1 gpc1_1_7970(
      {stage099[259]},
      {stage099[284]}
   );
   gpc1_1 gpc1_1_7971(
      {stage099[260]},
      {stage099[285]}
   );
   gpc1_1 gpc1_1_7972(
      {stage099[261]},
      {stage099[286]}
   );
   gpc606_5 gpc606_5_7973(
      {stage099[262], stage099[263], stage099[264], stage099[265], stage099[266], stage099[267]},
      {stage101[229], stage101[230], stage101[231], stage101[232], stage101[233], stage101[234]},
      {stage103[237], stage102[236], stage101[254], stage100[220], stage099[287]}
   );
   gpc606_5 gpc606_5_7974(
      {stage099[268], stage099[269], stage099[270], stage099[271], stage099[272], stage099[273]},
      {stage101[235], stage101[236], stage101[237], stage101[238], stage101[239], stage101[240]},
      {stage103[238], stage102[237], stage101[255], stage100[221], stage099[288]}
   );
   gpc606_5 gpc606_5_7975(
      {stage099[274], stage099[275], stage099[276], stage099[277], stage099[278], stage099[279]},
      {stage101[241], stage101[242], stage101[243], stage101[244], stage101[245], stage101[246]},
      {stage103[239], stage102[238], stage101[256], stage100[222], stage099[289]}
   );
   gpc606_5 gpc606_5_7976(
      {stage100[208], stage100[209], stage100[210], stage100[211], stage100[212], stage100[213]},
      {stage102[221], stage102[222], stage102[223], stage102[224], stage102[225], stage102[226]},
      {stage104[257], stage103[240], stage102[239], stage101[257], stage100[223]}
   );
   gpc606_5 gpc606_5_7977(
      {stage100[214], stage100[215], stage100[216], stage100[217], 1'h0, 1'h0},
      {stage102[227], stage102[228], stage102[229], stage102[230], stage102[231], stage102[232]},
      {stage104[258], stage103[241], stage102[240], stage101[258], stage100[224]}
   );
   gpc606_5 gpc606_5_7978(
      {stage101[247], stage101[248], stage101[249], stage101[250], stage101[251], stage101[252]},
      {stage103[225], stage103[226], stage103[227], stage103[228], stage103[229], stage103[230]},
      {stage105[217], stage104[259], stage103[242], stage102[241], stage101[259]}
   );
   gpc1_1 gpc1_1_7979(
      {stage102[233]},
      {stage102[242]}
   );
   gpc1_1 gpc1_1_7980(
      {stage102[234]},
      {stage102[243]}
   );
   gpc1_1 gpc1_1_7981(
      {stage103[231]},
      {stage103[243]}
   );
   gpc1_1 gpc1_1_7982(
      {stage103[232]},
      {stage103[244]}
   );
   gpc1_1 gpc1_1_7983(
      {stage103[233]},
      {stage103[245]}
   );
   gpc1_1 gpc1_1_7984(
      {stage103[234]},
      {stage103[246]}
   );
   gpc1_1 gpc1_1_7985(
      {stage103[235]},
      {stage103[247]}
   );
   gpc1_1 gpc1_1_7986(
      {stage103[236]},
      {stage103[248]}
   );
   gpc606_5 gpc606_5_7987(
      {stage104[245], stage104[246], stage104[247], stage104[248], stage104[249], stage104[250]},
      {stage106[229], stage106[230], stage106[231], stage106[232], stage106[233], stage106[234]},
      {stage108[247], stage107[248], stage106[248], stage105[218], stage104[260]}
   );
   gpc606_5 gpc606_5_7988(
      {stage104[251], stage104[252], stage104[253], stage104[254], stage104[255], stage104[256]},
      {stage106[235], stage106[236], stage106[237], stage106[238], stage106[239], stage106[240]},
      {stage108[248], stage107[249], stage106[249], stage105[219], stage104[261]}
   );
   gpc1_1 gpc1_1_7989(
      {stage105[206]},
      {stage105[220]}
   );
   gpc615_5 gpc615_5_7990(
      {stage105[207], stage105[208], stage105[209], stage105[210], stage105[211]},
      {stage106[241]},
      {stage107[228], stage107[229], stage107[230], stage107[231], stage107[232], stage107[233]},
      {stage109[224], stage108[249], stage107[250], stage106[250], stage105[221]}
   );
   gpc615_5 gpc615_5_7991(
      {stage105[212], stage105[213], stage105[214], stage105[215], stage105[216]},
      {stage106[242]},
      {stage107[234], stage107[235], stage107[236], stage107[237], stage107[238], stage107[239]},
      {stage109[225], stage108[250], stage107[251], stage106[251], stage105[222]}
   );
   gpc615_5 gpc615_5_7992(
      {stage106[243], stage106[244], stage106[245], stage106[246], stage106[247]},
      {stage107[240]},
      {stage108[225], stage108[226], stage108[227], stage108[228], stage108[229], stage108[230]},
      {stage110[256], stage109[226], stage108[251], stage107[252], stage106[252]}
   );
   gpc1_1 gpc1_1_7993(
      {stage107[241]},
      {stage107[253]}
   );
   gpc606_5 gpc606_5_7994(
      {stage107[242], stage107[243], stage107[244], stage107[245], stage107[246], stage107[247]},
      {stage109[209], stage109[210], stage109[211], stage109[212], stage109[213], stage109[214]},
      {stage111[254], stage110[257], stage109[227], stage108[252], stage107[254]}
   );
   gpc1_1 gpc1_1_7995(
      {stage108[231]},
      {stage108[253]}
   );
   gpc1_1 gpc1_1_7996(
      {stage108[232]},
      {stage108[254]}
   );
   gpc1_1 gpc1_1_7997(
      {stage108[233]},
      {stage108[255]}
   );
   gpc1_1 gpc1_1_7998(
      {stage108[234]},
      {stage108[256]}
   );
   gpc606_5 gpc606_5_7999(
      {stage108[235], stage108[236], stage108[237], stage108[238], stage108[239], stage108[240]},
      {stage110[236], stage110[237], stage110[238], stage110[239], stage110[240], stage110[241]},
      {stage112[227], stage111[255], stage110[258], stage109[228], stage108[257]}
   );
   gpc606_5 gpc606_5_8000(
      {stage108[241], stage108[242], stage108[243], stage108[244], stage108[245], stage108[246]},
      {stage110[242], stage110[243], stage110[244], stage110[245], stage110[246], stage110[247]},
      {stage112[228], stage111[256], stage110[259], stage109[229], stage108[258]}
   );
   gpc615_5 gpc615_5_8001(
      {stage109[215], stage109[216], stage109[217], stage109[218], stage109[219]},
      {stage110[248]},
      {stage111[242], stage111[243], stage111[244], stage111[245], stage111[246], stage111[247]},
      {stage113[226], stage112[229], stage111[257], stage110[260], stage109[230]}
   );
   gpc615_5 gpc615_5_8002(
      {stage109[220], stage109[221], stage109[222], stage109[223], 1'h0},
      {stage110[249]},
      {stage111[248], stage111[249], stage111[250], stage111[251], stage111[252], stage111[253]},
      {stage113[227], stage112[230], stage111[258], stage110[261], stage109[231]}
   );
   gpc1_1 gpc1_1_8003(
      {stage110[250]},
      {stage110[262]}
   );
   gpc1415_5 gpc1415_5_8004(
      {stage110[251], stage110[252], stage110[253], stage110[254], stage110[255]},
      {1'h0},
      {stage112[215], stage112[216], stage112[217], stage112[218]},
      {stage113[213]},
      {stage114[234], stage113[228], stage112[231], stage111[259], stage110[263]}
   );
   gpc1_1 gpc1_1_8005(
      {stage112[219]},
      {stage112[232]}
   );
   gpc1_1 gpc1_1_8006(
      {stage112[220]},
      {stage112[233]}
   );
   gpc606_5 gpc606_5_8007(
      {stage112[221], stage112[222], stage112[223], stage112[224], stage112[225], stage112[226]},
      {stage114[216], stage114[217], stage114[218], stage114[219], stage114[220], stage114[221]},
      {stage116[231], stage115[252], stage114[235], stage113[229], stage112[234]}
   );
   gpc1_1 gpc1_1_8008(
      {stage113[214]},
      {stage113[230]}
   );
   gpc1_1 gpc1_1_8009(
      {stage113[215]},
      {stage113[231]}
   );
   gpc1_1 gpc1_1_8010(
      {stage113[216]},
      {stage113[232]}
   );
   gpc1_1 gpc1_1_8011(
      {stage113[217]},
      {stage113[233]}
   );
   gpc1_1 gpc1_1_8012(
      {stage113[218]},
      {stage113[234]}
   );
   gpc1_1 gpc1_1_8013(
      {stage113[219]},
      {stage113[235]}
   );
   gpc606_5 gpc606_5_8014(
      {stage113[220], stage113[221], stage113[222], stage113[223], stage113[224], stage113[225]},
      {stage115[237], stage115[238], stage115[239], stage115[240], stage115[241], stage115[242]},
      {stage117[244], stage116[232], stage115[253], stage114[236], stage113[236]}
   );
   gpc606_5 gpc606_5_8015(
      {stage114[222], stage114[223], stage114[224], stage114[225], stage114[226], stage114[227]},
      {stage116[214], stage116[215], stage116[216], stage116[217], stage116[218], stage116[219]},
      {stage118[248], stage117[245], stage116[233], stage115[254], stage114[237]}
   );
   gpc606_5 gpc606_5_8016(
      {stage114[228], stage114[229], stage114[230], stage114[231], stage114[232], stage114[233]},
      {stage116[220], stage116[221], stage116[222], stage116[223], stage116[224], stage116[225]},
      {stage118[249], stage117[246], stage116[234], stage115[255], stage114[238]}
   );
   gpc623_5 gpc623_5_8017(
      {stage115[243], stage115[244], stage115[245]},
      {stage116[226], stage116[227]},
      {stage117[223], stage117[224], stage117[225], stage117[226], stage117[227], stage117[228]},
      {stage119[220], stage118[250], stage117[247], stage116[235], stage115[256]}
   );
   gpc623_5 gpc623_5_8018(
      {stage115[246], stage115[247], stage115[248]},
      {stage116[228], stage116[229]},
      {stage117[229], stage117[230], stage117[231], stage117[232], stage117[233], stage117[234]},
      {stage119[221], stage118[251], stage117[248], stage116[236], stage115[257]}
   );
   gpc623_5 gpc623_5_8019(
      {stage115[249], stage115[250], stage115[251]},
      {stage116[230], 1'h0},
      {stage117[235], stage117[236], stage117[237], stage117[238], stage117[239], stage117[240]},
      {stage119[222], stage118[252], stage117[249], stage116[237], stage115[258]}
   );
   gpc1_1 gpc1_1_8020(
      {stage117[241]},
      {stage117[250]}
   );
   gpc1_1 gpc1_1_8021(
      {stage117[242]},
      {stage117[251]}
   );
   gpc1_1 gpc1_1_8022(
      {stage117[243]},
      {stage117[252]}
   );
   gpc606_5 gpc606_5_8023(
      {stage118[224], stage118[225], stage118[226], stage118[227], stage118[228], stage118[229]},
      {stage120[220], stage120[221], stage120[222], stage120[223], stage120[224], stage120[225]},
      {stage122[235], stage121[217], stage120[245], stage119[223], stage118[253]}
   );
   gpc606_5 gpc606_5_8024(
      {stage118[230], stage118[231], stage118[232], stage118[233], stage118[234], stage118[235]},
      {stage120[226], stage120[227], stage120[228], stage120[229], stage120[230], stage120[231]},
      {stage122[236], stage121[218], stage120[246], stage119[224], stage118[254]}
   );
   gpc606_5 gpc606_5_8025(
      {stage118[236], stage118[237], stage118[238], stage118[239], stage118[240], stage118[241]},
      {stage120[232], stage120[233], stage120[234], stage120[235], stage120[236], stage120[237]},
      {stage122[237], stage121[219], stage120[247], stage119[225], stage118[255]}
   );
   gpc606_5 gpc606_5_8026(
      {stage118[242], stage118[243], stage118[244], stage118[245], stage118[246], stage118[247]},
      {stage120[238], stage120[239], stage120[240], stage120[241], stage120[242], stage120[243]},
      {stage122[238], stage121[220], stage120[248], stage119[226], stage118[256]}
   );
   gpc1_1 gpc1_1_8027(
      {stage119[210]},
      {stage119[227]}
   );
   gpc1_1 gpc1_1_8028(
      {stage119[211]},
      {stage119[228]}
   );
   gpc1_1 gpc1_1_8029(
      {stage119[212]},
      {stage119[229]}
   );
   gpc1_1 gpc1_1_8030(
      {stage119[213]},
      {stage119[230]}
   );
   gpc1406_5 gpc1406_5_8031(
      {stage119[214], stage119[215], stage119[216], stage119[217], stage119[218], stage119[219]},
      {stage121[205], stage121[206], stage121[207], stage121[208]},
      {stage122[222]},
      {stage123[306], stage122[239], stage121[221], stage120[249], stage119[231]}
   );
   gpc1_1 gpc1_1_8032(
      {stage120[244]},
      {stage120[250]}
   );
   gpc1_1 gpc1_1_8033(
      {stage121[209]},
      {stage121[222]}
   );
   gpc1_1 gpc1_1_8034(
      {stage121[210]},
      {stage121[223]}
   );
   gpc606_5 gpc606_5_8035(
      {stage121[211], stage121[212], stage121[213], stage121[214], stage121[215], stage121[216]},
      {stage123[282], stage123[283], stage123[284], stage123[285], stage123[286], stage123[287]},
      {stage125[263], stage124[224], stage123[307], stage122[240], stage121[224]}
   );
   gpc606_5 gpc606_5_8036(
      {stage122[223], stage122[224], stage122[225], stage122[226], stage122[227], stage122[228]},
      {stage124[212], stage124[213], stage124[214], stage124[215], stage124[216], stage124[217]},
      {stage126[263], stage125[264], stage124[225], stage123[308], stage122[241]}
   );
   gpc606_5 gpc606_5_8037(
      {stage122[229], stage122[230], stage122[231], stage122[232], stage122[233], stage122[234]},
      {stage124[218], stage124[219], stage124[220], stage124[221], stage124[222], stage124[223]},
      {stage126[264], stage125[265], stage124[226], stage123[309], stage122[242]}
   );
   gpc1_1 gpc1_1_8038(
      {stage123[288]},
      {stage123[310]}
   );
   gpc1_1 gpc1_1_8039(
      {stage123[289]},
      {stage123[311]}
   );
   gpc1_1 gpc1_1_8040(
      {stage123[290]},
      {stage123[312]}
   );
   gpc1_1 gpc1_1_8041(
      {stage123[291]},
      {stage123[313]}
   );
   gpc1_1 gpc1_1_8042(
      {stage123[292]},
      {stage123[314]}
   );
   gpc1_1 gpc1_1_8043(
      {stage123[293]},
      {stage123[315]}
   );
   gpc606_5 gpc606_5_8044(
      {stage123[294], stage123[295], stage123[296], stage123[297], stage123[298], stage123[299]},
      {stage125[241], stage125[242], stage125[243], stage125[244], stage125[245], stage125[246]},
      {stage127[268], stage126[265], stage125[266], stage124[227], stage123[316]}
   );
   gpc1406_5 gpc1406_5_8045(
      {stage123[300], stage123[301], stage123[302], stage123[303], stage123[304], stage123[305]},
      {stage125[247], stage125[248], stage125[249], stage125[250]},
      {stage126[242]},
      {stage127[269], stage126[266], stage125[267], stage124[228], stage123[317]}
   );
   gpc1_1 gpc1_1_8046(
      {stage125[251]},
      {stage125[268]}
   );
   gpc1_1 gpc1_1_8047(
      {stage125[252]},
      {stage125[269]}
   );
   gpc1_1 gpc1_1_8048(
      {stage125[253]},
      {stage125[270]}
   );
   gpc1_1 gpc1_1_8049(
      {stage125[254]},
      {stage125[271]}
   );
   gpc1_1 gpc1_1_8050(
      {stage125[255]},
      {stage125[272]}
   );
   gpc1_1 gpc1_1_8051(
      {stage125[256]},
      {stage125[273]}
   );
   gpc1_1 gpc1_1_8052(
      {stage125[257]},
      {stage125[274]}
   );
   gpc1_1 gpc1_1_8053(
      {stage125[258]},
      {stage125[275]}
   );
   gpc1_1 gpc1_1_8054(
      {stage125[259]},
      {stage125[276]}
   );
   gpc1_1 gpc1_1_8055(
      {stage125[260]},
      {stage125[277]}
   );
   gpc1_1 gpc1_1_8056(
      {stage125[261]},
      {stage125[278]}
   );
   gpc1_1 gpc1_1_8057(
      {stage125[262]},
      {stage125[279]}
   );
   gpc1_1 gpc1_1_8058(
      {stage126[243]},
      {stage126[267]}
   );
   gpc1_1 gpc1_1_8059(
      {stage126[244]},
      {stage126[268]}
   );
   gpc1_1 gpc1_1_8060(
      {stage126[245]},
      {stage126[269]}
   );
   gpc1_1 gpc1_1_8061(
      {stage126[246]},
      {stage126[270]}
   );
   gpc1_1 gpc1_1_8062(
      {stage126[247]},
      {stage126[271]}
   );
   gpc1_1 gpc1_1_8063(
      {stage126[248]},
      {stage126[272]}
   );
   gpc1_1 gpc1_1_8064(
      {stage126[249]},
      {stage126[273]}
   );
   gpc1_1 gpc1_1_8065(
      {stage126[250]},
      {stage126[274]}
   );
   gpc606_5 gpc606_5_8066(
      {stage126[251], stage126[252], stage126[253], stage126[254], stage126[255], stage126[256]},
      {stage128[47], stage128[48], stage128[49], stage128[50], stage128[51], stage128[52]},
      {stage130[9], stage129[56], stage128[72], stage127[270], stage126[275]}
   );
   gpc606_5 gpc606_5_8067(
      {stage126[257], stage126[258], stage126[259], stage126[260], stage126[261], stage126[262]},
      {stage128[53], stage128[54], stage128[55], stage128[56], stage128[57], stage128[58]},
      {stage130[10], stage129[57], stage128[73], stage127[271], stage126[276]}
   );
   gpc1_1 gpc1_1_8068(
      {stage127[254]},
      {stage127[272]}
   );
   gpc1_1 gpc1_1_8069(
      {stage127[255]},
      {stage127[273]}
   );
   gpc1_1 gpc1_1_8070(
      {stage127[256]},
      {stage127[274]}
   );
   gpc1_1 gpc1_1_8071(
      {stage127[257]},
      {stage127[275]}
   );
   gpc1_1 gpc1_1_8072(
      {stage127[258]},
      {stage127[276]}
   );
   gpc1_1 gpc1_1_8073(
      {stage127[259]},
      {stage127[277]}
   );
   gpc1_1 gpc1_1_8074(
      {stage127[260]},
      {stage127[278]}
   );
   gpc1_1 gpc1_1_8075(
      {stage127[261]},
      {stage127[279]}
   );
   gpc606_5 gpc606_5_8076(
      {stage127[262], stage127[263], stage127[264], stage127[265], stage127[266], stage127[267]},
      {stage129[39], stage129[40], stage129[41], stage129[42], stage129[43], stage129[44]},
      {stage131[4], stage130[11], stage129[58], stage128[74], stage127[280]}
   );
   gpc1_1 gpc1_1_8077(
      {stage128[59]},
      {stage128[75]}
   );
   gpc1_1 gpc1_1_8078(
      {stage128[60]},
      {stage128[76]}
   );
   gpc1_1 gpc1_1_8079(
      {stage128[61]},
      {stage128[77]}
   );
   gpc1_1 gpc1_1_8080(
      {stage128[62]},
      {stage128[78]}
   );
   gpc1_1 gpc1_1_8081(
      {stage128[63]},
      {stage128[79]}
   );
   gpc1_1 gpc1_1_8082(
      {stage128[64]},
      {stage128[80]}
   );
   gpc1_1 gpc1_1_8083(
      {stage128[65]},
      {stage128[81]}
   );
   gpc606_5 gpc606_5_8084(
      {stage128[66], stage128[67], stage128[68], stage128[69], stage128[70], stage128[71]},
      {stage130[5], stage130[6], stage130[7], stage130[8], 1'h0, 1'h0},
      {stage132[1], stage131[5], stage130[12], stage129[59], stage128[82]}
   );
   gpc1_1 gpc1_1_8085(
      {stage129[45]},
      {stage129[60]}
   );
   gpc1_1 gpc1_1_8086(
      {stage129[46]},
      {stage129[61]}
   );
   gpc1_1 gpc1_1_8087(
      {stage129[47]},
      {stage129[62]}
   );
   gpc1_1 gpc1_1_8088(
      {stage129[48]},
      {stage129[63]}
   );
   gpc1_1 gpc1_1_8089(
      {stage129[49]},
      {stage129[64]}
   );
   gpc606_5 gpc606_5_8090(
      {stage129[50], stage129[51], stage129[52], stage129[53], stage129[54], stage129[55]},
      {stage131[0], stage131[1], stage131[2], stage131[3], 1'h0, 1'h0},
      {stage133[0], stage132[2], stage131[6], stage130[13], stage129[65]}
   );
   gpc1_1 gpc1_1_8091(
      {stage132[0]},
      {stage132[3]}
   );
   gpc1_1 gpc1_1_8092(
      {stage000[186]},
      {stage000[188]}
   );
   gpc1_1 gpc1_1_8093(
      {stage000[187]},
      {stage000[189]}
   );
   gpc1_1 gpc1_1_8094(
      {stage001[218]},
      {stage001[226]}
   );
   gpc207_4 gpc207_4_8095(
      {stage001[219], stage001[220], stage001[221], stage001[222], stage001[223], stage001[224], stage001[225]},
      {stage003[206], stage003[207]},
      {stage004[263], stage003[214], stage002[242], stage001[227]}
   );
   gpc7_3 gpc7_3_8096(
      {stage002[235], stage002[236], stage002[237], stage002[238], stage002[239], stage002[240], stage002[241]},
      {stage004[264], stage003[215], stage002[243]}
   );
   gpc1343_5 gpc1343_5_8097(
      {stage003[208], stage003[209], stage003[210]},
      {stage004[252], stage004[253], stage004[254], stage004[255]},
      {stage005[263], stage005[264], stage005[265]},
      {stage006[245]},
      {stage007[250], stage006[251], stage005[277], stage004[265], stage003[216]}
   );
   gpc1343_5 gpc1343_5_8098(
      {stage003[211], stage003[212], stage003[213]},
      {stage004[256], stage004[257], stage004[258], stage004[259]},
      {stage005[266], stage005[267], stage005[268]},
      {stage006[246]},
      {stage007[251], stage006[252], stage005[278], stage004[266], stage003[217]}
   );
   gpc1_1 gpc1_1_8099(
      {stage004[260]},
      {stage004[267]}
   );
   gpc1_1 gpc1_1_8100(
      {stage004[261]},
      {stage004[268]}
   );
   gpc1_1 gpc1_1_8101(
      {stage004[262]},
      {stage004[269]}
   );
   gpc1_1 gpc1_1_8102(
      {stage005[269]},
      {stage005[279]}
   );
   gpc207_4 gpc207_4_8103(
      {stage005[270], stage005[271], stage005[272], stage005[273], stage005[274], stage005[275], stage005[276]},
      {stage007[244], stage007[245]},
      {stage008[236], stage007[252], stage006[253], stage005[280]}
   );
   gpc1_1 gpc1_1_8104(
      {stage006[247]},
      {stage006[254]}
   );
   gpc1_1 gpc1_1_8105(
      {stage006[248]},
      {stage006[255]}
   );
   gpc1_1 gpc1_1_8106(
      {stage006[249]},
      {stage006[256]}
   );
   gpc1_1 gpc1_1_8107(
      {stage006[250]},
      {stage006[257]}
   );
   gpc1_1 gpc1_1_8108(
      {stage007[246]},
      {stage007[253]}
   );
   gpc1_1 gpc1_1_8109(
      {stage007[247]},
      {stage007[254]}
   );
   gpc1_1 gpc1_1_8110(
      {stage007[248]},
      {stage007[255]}
   );
   gpc1_1 gpc1_1_8111(
      {stage007[249]},
      {stage007[256]}
   );
   gpc1_1 gpc1_1_8112(
      {stage008[223]},
      {stage008[237]}
   );
   gpc1_1 gpc1_1_8113(
      {stage008[224]},
      {stage008[238]}
   );
   gpc1_1 gpc1_1_8114(
      {stage008[225]},
      {stage008[239]}
   );
   gpc1_1 gpc1_1_8115(
      {stage008[226]},
      {stage008[240]}
   );
   gpc1_1 gpc1_1_8116(
      {stage008[227]},
      {stage008[241]}
   );
   gpc1_1 gpc1_1_8117(
      {stage008[228]},
      {stage008[242]}
   );
   gpc1_1 gpc1_1_8118(
      {stage008[229]},
      {stage008[243]}
   );
   gpc606_5 gpc606_5_8119(
      {stage008[230], stage008[231], stage008[232], stage008[233], stage008[234], stage008[235]},
      {stage010[279], stage010[280], stage010[281], stage010[282], stage010[283], stage010[284]},
      {stage012[319], stage011[254], stage010[291], stage009[237], stage008[244]}
   );
   gpc606_5 gpc606_5_8120(
      {stage009[231], stage009[232], stage009[233], stage009[234], stage009[235], stage009[236]},
      {stage011[239], stage011[240], stage011[241], stage011[242], stage011[243], stage011[244]},
      {stage013[253], stage012[320], stage011[255], stage010[292], stage009[238]}
   );
   gpc1_1 gpc1_1_8121(
      {stage010[285]},
      {stage010[293]}
   );
   gpc1_1 gpc1_1_8122(
      {stage010[286]},
      {stage010[294]}
   );
   gpc1_1 gpc1_1_8123(
      {stage010[287]},
      {stage010[295]}
   );
   gpc1_1 gpc1_1_8124(
      {stage010[288]},
      {stage010[296]}
   );
   gpc1_1 gpc1_1_8125(
      {stage010[289]},
      {stage010[297]}
   );
   gpc1_1 gpc1_1_8126(
      {stage010[290]},
      {stage010[298]}
   );
   gpc1_1 gpc1_1_8127(
      {stage011[245]},
      {stage011[256]}
   );
   gpc1_1 gpc1_1_8128(
      {stage011[246]},
      {stage011[257]}
   );
   gpc1_1 gpc1_1_8129(
      {stage011[247]},
      {stage011[258]}
   );
   gpc1_1 gpc1_1_8130(
      {stage011[248]},
      {stage011[259]}
   );
   gpc615_5 gpc615_5_8131(
      {stage011[249], stage011[250], stage011[251], stage011[252], stage011[253]},
      {stage012[310]},
      {stage013[235], stage013[236], stage013[237], stage013[238], stage013[239], stage013[240]},
      {stage015[253], stage014[298], stage013[254], stage012[321], stage011[260]}
   );
   gpc1_1 gpc1_1_8132(
      {stage012[311]},
      {stage012[322]}
   );
   gpc1_1 gpc1_1_8133(
      {stage012[312]},
      {stage012[323]}
   );
   gpc606_5 gpc606_5_8134(
      {stage012[313], stage012[314], stage012[315], stage012[316], stage012[317], stage012[318]},
      {stage014[288], stage014[289], stage014[290], stage014[291], stage014[292], stage014[293]},
      {stage016[285], stage015[254], stage014[299], stage013[255], stage012[324]}
   );
   gpc1_1 gpc1_1_8135(
      {stage013[241]},
      {stage013[256]}
   );
   gpc1_1 gpc1_1_8136(
      {stage013[242]},
      {stage013[257]}
   );
   gpc1_1 gpc1_1_8137(
      {stage013[243]},
      {stage013[258]}
   );
   gpc1_1 gpc1_1_8138(
      {stage013[244]},
      {stage013[259]}
   );
   gpc1_1 gpc1_1_8139(
      {stage013[245]},
      {stage013[260]}
   );
   gpc1_1 gpc1_1_8140(
      {stage013[246]},
      {stage013[261]}
   );
   gpc1_1 gpc1_1_8141(
      {stage013[247]},
      {stage013[262]}
   );
   gpc1_1 gpc1_1_8142(
      {stage013[248]},
      {stage013[263]}
   );
   gpc1_1 gpc1_1_8143(
      {stage013[249]},
      {stage013[264]}
   );
   gpc1_1 gpc1_1_8144(
      {stage013[250]},
      {stage013[265]}
   );
   gpc1_1 gpc1_1_8145(
      {stage013[251]},
      {stage013[266]}
   );
   gpc1_1 gpc1_1_8146(
      {stage013[252]},
      {stage013[267]}
   );
   gpc1_1 gpc1_1_8147(
      {stage014[294]},
      {stage014[300]}
   );
   gpc1_1 gpc1_1_8148(
      {stage014[295]},
      {stage014[301]}
   );
   gpc1_1 gpc1_1_8149(
      {stage014[296]},
      {stage014[302]}
   );
   gpc1_1 gpc1_1_8150(
      {stage014[297]},
      {stage014[303]}
   );
   gpc1_1 gpc1_1_8151(
      {stage015[240]},
      {stage015[255]}
   );
   gpc1_1 gpc1_1_8152(
      {stage015[241]},
      {stage015[256]}
   );
   gpc1_1 gpc1_1_8153(
      {stage015[242]},
      {stage015[257]}
   );
   gpc615_5 gpc615_5_8154(
      {stage015[243], stage015[244], stage015[245], stage015[246], stage015[247]},
      {stage016[275]},
      {stage017[266], stage017[267], stage017[268], stage017[269], stage017[270], stage017[271]},
      {stage019[258], stage018[249], stage017[278], stage016[286], stage015[258]}
   );
   gpc615_5 gpc615_5_8155(
      {stage015[248], stage015[249], stage015[250], stage015[251], stage015[252]},
      {stage016[276]},
      {stage017[272], stage017[273], stage017[274], stage017[275], stage017[276], stage017[277]},
      {stage019[259], stage018[250], stage017[279], stage016[287], stage015[259]}
   );
   gpc1_1 gpc1_1_8156(
      {stage016[277]},
      {stage016[288]}
   );
   gpc1_1 gpc1_1_8157(
      {stage016[278]},
      {stage016[289]}
   );
   gpc606_5 gpc606_5_8158(
      {stage016[279], stage016[280], stage016[281], stage016[282], stage016[283], stage016[284]},
      {stage018[241], stage018[242], stage018[243], stage018[244], stage018[245], stage018[246]},
      {stage020[229], stage019[260], stage018[251], stage017[280], stage016[290]}
   );
   gpc1_1 gpc1_1_8159(
      {stage018[247]},
      {stage018[252]}
   );
   gpc1_1 gpc1_1_8160(
      {stage018[248]},
      {stage018[253]}
   );
   gpc1_1 gpc1_1_8161(
      {stage019[246]},
      {stage019[261]}
   );
   gpc1_1 gpc1_1_8162(
      {stage019[247]},
      {stage019[262]}
   );
   gpc1_1 gpc1_1_8163(
      {stage019[248]},
      {stage019[263]}
   );
   gpc1_1 gpc1_1_8164(
      {stage019[249]},
      {stage019[264]}
   );
   gpc1_1 gpc1_1_8165(
      {stage019[250]},
      {stage019[265]}
   );
   gpc1_1 gpc1_1_8166(
      {stage019[251]},
      {stage019[266]}
   );
   gpc1_1 gpc1_1_8167(
      {stage019[252]},
      {stage019[267]}
   );
   gpc615_5 gpc615_5_8168(
      {stage019[253], stage019[254], stage019[255], stage019[256], stage019[257]},
      {stage020[219]},
      {stage021[271], stage021[272], stage021[273], stage021[274], stage021[275], stage021[276]},
      {stage023[309], stage022[225], stage021[285], stage020[230], stage019[268]}
   );
   gpc1_1 gpc1_1_8169(
      {stage020[220]},
      {stage020[231]}
   );
   gpc1_1 gpc1_1_8170(
      {stage020[221]},
      {stage020[232]}
   );
   gpc1_1 gpc1_1_8171(
      {stage020[222]},
      {stage020[233]}
   );
   gpc606_5 gpc606_5_8172(
      {stage020[223], stage020[224], stage020[225], stage020[226], stage020[227], stage020[228]},
      {stage022[215], stage022[216], stage022[217], stage022[218], stage022[219], stage022[220]},
      {stage024[254], stage023[310], stage022[226], stage021[286], stage020[234]}
   );
   gpc1_1 gpc1_1_8173(
      {stage021[277]},
      {stage021[287]}
   );
   gpc1_1 gpc1_1_8174(
      {stage021[278]},
      {stage021[288]}
   );
   gpc1_1 gpc1_1_8175(
      {stage021[279]},
      {stage021[289]}
   );
   gpc1_1 gpc1_1_8176(
      {stage021[280]},
      {stage021[290]}
   );
   gpc1_1 gpc1_1_8177(
      {stage021[281]},
      {stage021[291]}
   );
   gpc1_1 gpc1_1_8178(
      {stage021[282]},
      {stage021[292]}
   );
   gpc1_1 gpc1_1_8179(
      {stage021[283]},
      {stage021[293]}
   );
   gpc1_1 gpc1_1_8180(
      {stage021[284]},
      {stage021[294]}
   );
   gpc1_1 gpc1_1_8181(
      {stage022[221]},
      {stage022[227]}
   );
   gpc1_1 gpc1_1_8182(
      {stage022[222]},
      {stage022[228]}
   );
   gpc1_1 gpc1_1_8183(
      {stage022[223]},
      {stage022[229]}
   );
   gpc1_1 gpc1_1_8184(
      {stage022[224]},
      {stage022[230]}
   );
   gpc1_1 gpc1_1_8185(
      {stage023[295]},
      {stage023[311]}
   );
   gpc1_1 gpc1_1_8186(
      {stage023[296]},
      {stage023[312]}
   );
   gpc1_1 gpc1_1_8187(
      {stage023[297]},
      {stage023[313]}
   );
   gpc1_1 gpc1_1_8188(
      {stage023[298]},
      {stage023[314]}
   );
   gpc615_5 gpc615_5_8189(
      {stage023[299], stage023[300], stage023[301], stage023[302], stage023[303]},
      {stage024[245]},
      {stage025[279], stage025[280], stage025[281], stage025[282], stage025[283], stage025[284]},
      {stage027[235], stage026[240], stage025[292], stage024[255], stage023[315]}
   );
   gpc615_5 gpc615_5_8190(
      {stage023[304], stage023[305], stage023[306], stage023[307], stage023[308]},
      {stage024[246]},
      {stage025[285], stage025[286], stage025[287], stage025[288], stage025[289], stage025[290]},
      {stage027[236], stage026[241], stage025[293], stage024[256], stage023[316]}
   );
   gpc1_1 gpc1_1_8191(
      {stage024[247]},
      {stage024[257]}
   );
   gpc606_5 gpc606_5_8192(
      {stage024[248], stage024[249], stage024[250], stage024[251], stage024[252], stage024[253]},
      {stage026[234], stage026[235], stage026[236], stage026[237], stage026[238], stage026[239]},
      {stage028[254], stage027[237], stage026[242], stage025[294], stage024[258]}
   );
   gpc1_1 gpc1_1_8193(
      {stage025[291]},
      {stage025[295]}
   );
   gpc1_1 gpc1_1_8194(
      {stage027[229]},
      {stage027[238]}
   );
   gpc615_5 gpc615_5_8195(
      {stage027[230], stage027[231], stage027[232], stage027[233], stage027[234]},
      {stage028[239]},
      {stage029[274], stage029[275], stage029[276], stage029[277], stage029[278], stage029[279]},
      {stage031[250], stage030[240], stage029[285], stage028[255], stage027[239]}
   );
   gpc1_1 gpc1_1_8196(
      {stage028[240]},
      {stage028[256]}
   );
   gpc1_1 gpc1_1_8197(
      {stage028[241]},
      {stage028[257]}
   );
   gpc1_1 gpc1_1_8198(
      {stage028[242]},
      {stage028[258]}
   );
   gpc1_1 gpc1_1_8199(
      {stage028[243]},
      {stage028[259]}
   );
   gpc1_1 gpc1_1_8200(
      {stage028[244]},
      {stage028[260]}
   );
   gpc1_1 gpc1_1_8201(
      {stage028[245]},
      {stage028[261]}
   );
   gpc1_1 gpc1_1_8202(
      {stage028[246]},
      {stage028[262]}
   );
   gpc1_1 gpc1_1_8203(
      {stage028[247]},
      {stage028[263]}
   );
   gpc606_5 gpc606_5_8204(
      {stage028[248], stage028[249], stage028[250], stage028[251], stage028[252], stage028[253]},
      {stage030[230], stage030[231], stage030[232], stage030[233], stage030[234], stage030[235]},
      {stage032[298], stage031[251], stage030[241], stage029[286], stage028[264]}
   );
   gpc606_5 gpc606_5_8205(
      {stage029[280], stage029[281], stage029[282], stage029[283], stage029[284], 1'h0},
      {stage031[238], stage031[239], stage031[240], stage031[241], stage031[242], stage031[243]},
      {stage033[291], stage032[299], stage031[252], stage030[242], stage029[287]}
   );
   gpc1_1 gpc1_1_8206(
      {stage030[236]},
      {stage030[243]}
   );
   gpc1_1 gpc1_1_8207(
      {stage030[237]},
      {stage030[244]}
   );
   gpc1_1 gpc1_1_8208(
      {stage030[238]},
      {stage030[245]}
   );
   gpc1_1 gpc1_1_8209(
      {stage030[239]},
      {stage030[246]}
   );
   gpc1_1 gpc1_1_8210(
      {stage031[244]},
      {stage031[253]}
   );
   gpc615_5 gpc615_5_8211(
      {stage031[245], stage031[246], stage031[247], stage031[248], stage031[249]},
      {stage032[284]},
      {stage033[284], stage033[285], stage033[286], stage033[287], stage033[288], stage033[289]},
      {stage035[260], stage034[299], stage033[292], stage032[300], stage031[254]}
   );
   gpc1_1 gpc1_1_8212(
      {stage032[285]},
      {stage032[301]}
   );
   gpc606_5 gpc606_5_8213(
      {stage032[286], stage032[287], stage032[288], stage032[289], stage032[290], stage032[291]},
      {stage034[280], stage034[281], stage034[282], stage034[283], stage034[284], stage034[285]},
      {stage036[225], stage035[261], stage034[300], stage033[293], stage032[302]}
   );
   gpc606_5 gpc606_5_8214(
      {stage032[292], stage032[293], stage032[294], stage032[295], stage032[296], stage032[297]},
      {stage034[286], stage034[287], stage034[288], stage034[289], stage034[290], stage034[291]},
      {stage036[226], stage035[262], stage034[301], stage033[294], stage032[303]}
   );
   gpc1_1 gpc1_1_8215(
      {stage033[290]},
      {stage033[295]}
   );
   gpc1_1 gpc1_1_8216(
      {stage034[292]},
      {stage034[302]}
   );
   gpc1_1 gpc1_1_8217(
      {stage034[293]},
      {stage034[303]}
   );
   gpc1_1 gpc1_1_8218(
      {stage034[294]},
      {stage034[304]}
   );
   gpc1_1 gpc1_1_8219(
      {stage034[295]},
      {stage034[305]}
   );
   gpc1_1 gpc1_1_8220(
      {stage034[296]},
      {stage034[306]}
   );
   gpc1_1 gpc1_1_8221(
      {stage034[297]},
      {stage034[307]}
   );
   gpc1_1 gpc1_1_8222(
      {stage034[298]},
      {stage034[308]}
   );
   gpc1_1 gpc1_1_8223(
      {stage035[254]},
      {stage035[263]}
   );
   gpc615_5 gpc615_5_8224(
      {stage035[255], stage035[256], stage035[257], stage035[258], stage035[259]},
      {stage036[216]},
      {stage037[259], stage037[260], stage037[261], stage037[262], stage037[263], stage037[264]},
      {stage039[250], stage038[250], stage037[271], stage036[227], stage035[264]}
   );
   gpc1_1 gpc1_1_8225(
      {stage036[217]},
      {stage036[228]}
   );
   gpc1_1 gpc1_1_8226(
      {stage036[218]},
      {stage036[229]}
   );
   gpc606_5 gpc606_5_8227(
      {stage036[219], stage036[220], stage036[221], stage036[222], stage036[223], stage036[224]},
      {stage038[234], stage038[235], stage038[236], stage038[237], stage038[238], stage038[239]},
      {stage040[301], stage039[251], stage038[251], stage037[272], stage036[230]}
   );
   gpc1_1 gpc1_1_8228(
      {stage037[265]},
      {stage037[273]}
   );
   gpc1_1 gpc1_1_8229(
      {stage037[266]},
      {stage037[274]}
   );
   gpc1_1 gpc1_1_8230(
      {stage037[267]},
      {stage037[275]}
   );
   gpc1_1 gpc1_1_8231(
      {stage037[268]},
      {stage037[276]}
   );
   gpc1_1 gpc1_1_8232(
      {stage037[269]},
      {stage037[277]}
   );
   gpc1_1 gpc1_1_8233(
      {stage037[270]},
      {stage037[278]}
   );
   gpc1_1 gpc1_1_8234(
      {stage038[240]},
      {stage038[252]}
   );
   gpc1_1 gpc1_1_8235(
      {stage038[241]},
      {stage038[253]}
   );
   gpc1_1 gpc1_1_8236(
      {stage038[242]},
      {stage038[254]}
   );
   gpc1_1 gpc1_1_8237(
      {stage038[243]},
      {stage038[255]}
   );
   gpc606_5 gpc606_5_8238(
      {stage038[244], stage038[245], stage038[246], stage038[247], stage038[248], stage038[249]},
      {stage040[286], stage040[287], stage040[288], stage040[289], stage040[290], stage040[291]},
      {stage042[291], stage041[267], stage040[302], stage039[252], stage038[256]}
   );
   gpc1_1 gpc1_1_8239(
      {stage039[243]},
      {stage039[253]}
   );
   gpc1_1 gpc1_1_8240(
      {stage039[244]},
      {stage039[254]}
   );
   gpc615_5 gpc615_5_8241(
      {stage039[245], stage039[246], stage039[247], stage039[248], stage039[249]},
      {stage040[292]},
      {stage041[253], stage041[254], stage041[255], stage041[256], stage041[257], stage041[258]},
      {stage043[217], stage042[292], stage041[268], stage040[303], stage039[255]}
   );
   gpc1_1 gpc1_1_8242(
      {stage040[293]},
      {stage040[304]}
   );
   gpc1_1 gpc1_1_8243(
      {stage040[294]},
      {stage040[305]}
   );
   gpc606_5 gpc606_5_8244(
      {stage040[295], stage040[296], stage040[297], stage040[298], stage040[299], stage040[300]},
      {stage042[279], stage042[280], stage042[281], stage042[282], stage042[283], stage042[284]},
      {stage044[226], stage043[218], stage042[293], stage041[269], stage040[306]}
   );
   gpc1_1 gpc1_1_8245(
      {stage041[259]},
      {stage041[270]}
   );
   gpc1_1 gpc1_1_8246(
      {stage041[260]},
      {stage041[271]}
   );
   gpc1_1 gpc1_1_8247(
      {stage041[261]},
      {stage041[272]}
   );
   gpc1_1 gpc1_1_8248(
      {stage041[262]},
      {stage041[273]}
   );
   gpc1_1 gpc1_1_8249(
      {stage041[263]},
      {stage041[274]}
   );
   gpc1_1 gpc1_1_8250(
      {stage041[264]},
      {stage041[275]}
   );
   gpc1_1 gpc1_1_8251(
      {stage041[265]},
      {stage041[276]}
   );
   gpc1_1 gpc1_1_8252(
      {stage041[266]},
      {stage041[277]}
   );
   gpc1_1 gpc1_1_8253(
      {stage042[285]},
      {stage042[294]}
   );
   gpc615_5 gpc615_5_8254(
      {stage042[286], stage042[287], stage042[288], stage042[289], stage042[290]},
      {stage043[210]},
      {stage044[220], stage044[221], stage044[222], stage044[223], stage044[224], stage044[225]},
      {stage046[272], stage045[272], stage044[227], stage043[219], stage042[295]}
   );
   gpc606_5 gpc606_5_8255(
      {stage043[211], stage043[212], stage043[213], stage043[214], stage043[215], stage043[216]},
      {stage045[266], stage045[267], stage045[268], stage045[269], stage045[270], stage045[271]},
      {stage047[232], stage046[273], stage045[273], stage044[228], stage043[220]}
   );
   gpc1_1 gpc1_1_8256(
      {stage046[263]},
      {stage046[274]}
   );
   gpc1_1 gpc1_1_8257(
      {stage046[264]},
      {stage046[275]}
   );
   gpc1_1 gpc1_1_8258(
      {stage046[265]},
      {stage046[276]}
   );
   gpc1_1 gpc1_1_8259(
      {stage046[266]},
      {stage046[277]}
   );
   gpc615_5 gpc615_5_8260(
      {stage046[267], stage046[268], stage046[269], stage046[270], stage046[271]},
      {stage047[224]},
      {stage048[321], stage048[322], stage048[323], stage048[324], stage048[325], stage048[326]},
      {stage050[278], stage049[255], stage048[336], stage047[233], stage046[278]}
   );
   gpc1_1 gpc1_1_8261(
      {stage047[225]},
      {stage047[234]}
   );
   gpc1_1 gpc1_1_8262(
      {stage047[226]},
      {stage047[235]}
   );
   gpc615_5 gpc615_5_8263(
      {stage047[227], stage047[228], stage047[229], stage047[230], stage047[231]},
      {stage048[327]},
      {stage049[245], stage049[246], stage049[247], stage049[248], stage049[249], stage049[250]},
      {stage051[249], stage050[279], stage049[256], stage048[337], stage047[236]}
   );
   gpc1_1 gpc1_1_8264(
      {stage048[328]},
      {stage048[338]}
   );
   gpc1_1 gpc1_1_8265(
      {stage048[329]},
      {stage048[339]}
   );
   gpc1_1 gpc1_1_8266(
      {stage048[330]},
      {stage048[340]}
   );
   gpc1_1 gpc1_1_8267(
      {stage048[331]},
      {stage048[341]}
   );
   gpc1_1 gpc1_1_8268(
      {stage048[332]},
      {stage048[342]}
   );
   gpc1_1 gpc1_1_8269(
      {stage048[333]},
      {stage048[343]}
   );
   gpc1_1 gpc1_1_8270(
      {stage048[334]},
      {stage048[344]}
   );
   gpc1_1 gpc1_1_8271(
      {stage048[335]},
      {stage048[345]}
   );
   gpc615_5 gpc615_5_8272(
      {stage049[251], stage049[252], stage049[253], stage049[254], 1'h0},
      {stage050[268]},
      {stage051[237], stage051[238], stage051[239], stage051[240], stage051[241], stage051[242]},
      {stage053[249], stage052[274], stage051[250], stage050[280], stage049[257]}
   );
   gpc615_5 gpc615_5_8273(
      {stage050[269], stage050[270], stage050[271], stage050[272], stage050[273]},
      {stage051[243]},
      {stage052[263], stage052[264], stage052[265], stage052[266], stage052[267], stage052[268]},
      {stage054[255], stage053[250], stage052[275], stage051[251], stage050[281]}
   );
   gpc615_5 gpc615_5_8274(
      {stage050[274], stage050[275], stage050[276], stage050[277], 1'h0},
      {stage051[244]},
      {stage052[269], stage052[270], stage052[271], stage052[272], stage052[273], 1'h0},
      {stage054[256], stage053[251], stage052[276], stage051[252], stage050[282]}
   );
   gpc615_5 gpc615_5_8275(
      {stage051[245], stage051[246], stage051[247], stage051[248], 1'h0},
      {1'h0},
      {stage053[232], stage053[233], stage053[234], stage053[235], stage053[236], stage053[237]},
      {stage055[284], stage054[257], stage053[252], stage052[277], stage051[253]}
   );
   gpc606_5 gpc606_5_8276(
      {stage053[238], stage053[239], stage053[240], stage053[241], stage053[242], stage053[243]},
      {stage055[265], stage055[266], stage055[267], stage055[268], stage055[269], stage055[270]},
      {stage057[252], stage056[286], stage055[285], stage054[258], stage053[253]}
   );
   gpc606_5 gpc606_5_8277(
      {stage053[244], stage053[245], stage053[246], stage053[247], stage053[248], 1'h0},
      {stage055[271], stage055[272], stage055[273], stage055[274], stage055[275], stage055[276]},
      {stage057[253], stage056[287], stage055[286], stage054[259], stage053[254]}
   );
   gpc606_5 gpc606_5_8278(
      {stage054[245], stage054[246], stage054[247], stage054[248], stage054[249], stage054[250]},
      {stage056[263], stage056[264], stage056[265], stage056[266], stage056[267], stage056[268]},
      {stage058[232], stage057[254], stage056[288], stage055[287], stage054[260]}
   );
   gpc615_5 gpc615_5_8279(
      {stage054[251], stage054[252], stage054[253], stage054[254], 1'h0},
      {stage055[277]},
      {stage056[269], stage056[270], stage056[271], stage056[272], stage056[273], stage056[274]},
      {stage058[233], stage057[255], stage056[289], stage055[288], stage054[261]}
   );
   gpc1_1 gpc1_1_8280(
      {stage055[278]},
      {stage055[289]}
   );
   gpc1_1 gpc1_1_8281(
      {stage055[279]},
      {stage055[290]}
   );
   gpc1_1 gpc1_1_8282(
      {stage055[280]},
      {stage055[291]}
   );
   gpc1_1 gpc1_1_8283(
      {stage055[281]},
      {stage055[292]}
   );
   gpc1_1 gpc1_1_8284(
      {stage055[282]},
      {stage055[293]}
   );
   gpc1_1 gpc1_1_8285(
      {stage055[283]},
      {stage055[294]}
   );
   gpc606_5 gpc606_5_8286(
      {stage056[275], stage056[276], stage056[277], stage056[278], stage056[279], stage056[280]},
      {stage058[222], stage058[223], stage058[224], stage058[225], stage058[226], stage058[227]},
      {stage060[240], stage059[313], stage058[234], stage057[256], stage056[290]}
   );
   gpc606_5 gpc606_5_8287(
      {stage056[281], stage056[282], stage056[283], stage056[284], stage056[285], 1'h0},
      {stage058[228], stage058[229], stage058[230], stage058[231], 1'h0, 1'h0},
      {stage060[241], stage059[314], stage058[235], stage057[257], stage056[291]}
   );
   gpc606_5 gpc606_5_8288(
      {stage057[246], stage057[247], stage057[248], stage057[249], stage057[250], stage057[251]},
      {stage059[297], stage059[298], stage059[299], stage059[300], stage059[301], stage059[302]},
      {stage061[276], stage060[242], stage059[315], stage058[236], stage057[258]}
   );
   gpc1_1 gpc1_1_8289(
      {stage059[303]},
      {stage059[316]}
   );
   gpc1_1 gpc1_1_8290(
      {stage059[304]},
      {stage059[317]}
   );
   gpc1_1 gpc1_1_8291(
      {stage059[305]},
      {stage059[318]}
   );
   gpc1_1 gpc1_1_8292(
      {stage059[306]},
      {stage059[319]}
   );
   gpc606_5 gpc606_5_8293(
      {stage059[307], stage059[308], stage059[309], stage059[310], stage059[311], stage059[312]},
      {stage061[262], stage061[263], stage061[264], stage061[265], stage061[266], stage061[267]},
      {stage063[215], stage062[253], stage061[277], stage060[243], stage059[320]}
   );
   gpc1_1 gpc1_1_8294(
      {stage060[229]},
      {stage060[244]}
   );
   gpc615_5 gpc615_5_8295(
      {stage060[230], stage060[231], stage060[232], stage060[233], stage060[234]},
      {stage061[268]},
      {stage062[239], stage062[240], stage062[241], stage062[242], stage062[243], stage062[244]},
      {stage064[264], stage063[216], stage062[254], stage061[278], stage060[245]}
   );
   gpc615_5 gpc615_5_8296(
      {stage060[235], stage060[236], stage060[237], stage060[238], stage060[239]},
      {stage061[269]},
      {stage062[245], stage062[246], stage062[247], stage062[248], stage062[249], stage062[250]},
      {stage064[265], stage063[217], stage062[255], stage061[279], stage060[246]}
   );
   gpc606_5 gpc606_5_8297(
      {stage061[270], stage061[271], stage061[272], stage061[273], stage061[274], stage061[275]},
      {stage063[209], stage063[210], stage063[211], stage063[212], stage063[213], stage063[214]},
      {stage065[261], stage064[266], stage063[218], stage062[256], stage061[280]}
   );
   gpc1_1 gpc1_1_8298(
      {stage062[251]},
      {stage062[257]}
   );
   gpc1_1 gpc1_1_8299(
      {stage062[252]},
      {stage062[258]}
   );
   gpc1_1 gpc1_1_8300(
      {stage064[257]},
      {stage064[267]}
   );
   gpc606_5 gpc606_5_8301(
      {stage064[258], stage064[259], stage064[260], stage064[261], stage064[262], stage064[263]},
      {stage066[273], stage066[274], stage066[275], stage066[276], stage066[277], stage066[278]},
      {stage068[277], stage067[262], stage066[286], stage065[262], stage064[268]}
   );
   gpc606_5 gpc606_5_8302(
      {stage065[255], stage065[256], stage065[257], stage065[258], stage065[259], stage065[260]},
      {stage067[253], stage067[254], stage067[255], stage067[256], stage067[257], stage067[258]},
      {stage069[263], stage068[278], stage067[263], stage066[287], stage065[263]}
   );
   gpc1_1 gpc1_1_8303(
      {stage066[279]},
      {stage066[288]}
   );
   gpc606_5 gpc606_5_8304(
      {stage066[280], stage066[281], stage066[282], stage066[283], stage066[284], stage066[285]},
      {stage068[266], stage068[267], stage068[268], stage068[269], stage068[270], stage068[271]},
      {stage070[259], stage069[264], stage068[279], stage067[264], stage066[289]}
   );
   gpc1_1 gpc1_1_8305(
      {stage067[259]},
      {stage067[265]}
   );
   gpc1_1 gpc1_1_8306(
      {stage067[260]},
      {stage067[266]}
   );
   gpc1_1 gpc1_1_8307(
      {stage067[261]},
      {stage067[267]}
   );
   gpc615_5 gpc615_5_8308(
      {stage068[272], stage068[273], stage068[274], stage068[275], stage068[276]},
      {stage069[256]},
      {stage070[249], stage070[250], stage070[251], stage070[252], stage070[253], stage070[254]},
      {stage072[311], stage071[263], stage070[260], stage069[265], stage068[280]}
   );
   gpc1_1 gpc1_1_8309(
      {stage069[257]},
      {stage069[266]}
   );
   gpc1_1 gpc1_1_8310(
      {stage069[258]},
      {stage069[267]}
   );
   gpc1_1 gpc1_1_8311(
      {stage069[259]},
      {stage069[268]}
   );
   gpc1_1 gpc1_1_8312(
      {stage069[260]},
      {stage069[269]}
   );
   gpc1_1 gpc1_1_8313(
      {stage069[261]},
      {stage069[270]}
   );
   gpc1_1 gpc1_1_8314(
      {stage069[262]},
      {stage069[271]}
   );
   gpc1_1 gpc1_1_8315(
      {stage070[255]},
      {stage070[261]}
   );
   gpc1_1 gpc1_1_8316(
      {stage070[256]},
      {stage070[262]}
   );
   gpc1_1 gpc1_1_8317(
      {stage070[257]},
      {stage070[263]}
   );
   gpc1_1 gpc1_1_8318(
      {stage070[258]},
      {stage070[264]}
   );
   gpc1_1 gpc1_1_8319(
      {stage071[256]},
      {stage071[264]}
   );
   gpc606_5 gpc606_5_8320(
      {stage071[257], stage071[258], stage071[259], stage071[260], stage071[261], stage071[262]},
      {stage073[232], stage073[233], stage073[234], stage073[235], stage073[236], stage073[237]},
      {stage075[209], stage074[254], stage073[243], stage072[312], stage071[265]}
   );
   gpc7_3 gpc7_3_8321(
      {stage072[299], stage072[300], stage072[301], stage072[302], stage072[303], stage072[304], stage072[305]},
      {stage074[255], stage073[244], stage072[313]}
   );
   gpc606_5 gpc606_5_8322(
      {stage072[306], stage072[307], stage072[308], stage072[309], stage072[310], 1'h0},
      {stage074[243], stage074[244], stage074[245], stage074[246], stage074[247], stage074[248]},
      {stage076[215], stage075[210], stage074[256], stage073[245], stage072[314]}
   );
   gpc615_5 gpc615_5_8323(
      {stage073[238], stage073[239], stage073[240], stage073[241], stage073[242]},
      {stage074[249]},
      {stage075[205], stage075[206], stage075[207], stage075[208], 1'h0, 1'h0},
      {stage077[252], stage076[216], stage075[211], stage074[257], stage073[246]}
   );
   gpc1_1 gpc1_1_8324(
      {stage074[250]},
      {stage074[258]}
   );
   gpc1_1 gpc1_1_8325(
      {stage074[251]},
      {stage074[259]}
   );
   gpc1_1 gpc1_1_8326(
      {stage074[252]},
      {stage074[260]}
   );
   gpc1_1 gpc1_1_8327(
      {stage074[253]},
      {stage074[261]}
   );
   gpc606_5 gpc606_5_8328(
      {stage076[209], stage076[210], stage076[211], stage076[212], stage076[213], stage076[214]},
      {stage078[228], stage078[229], stage078[230], stage078[231], stage078[232], stage078[233]},
      {stage080[261], stage079[253], stage078[234], stage077[253], stage076[217]}
   );
   gpc1_1 gpc1_1_8329(
      {stage077[243]},
      {stage077[254]}
   );
   gpc1_1 gpc1_1_8330(
      {stage077[244]},
      {stage077[255]}
   );
   gpc1_1 gpc1_1_8331(
      {stage077[245]},
      {stage077[256]}
   );
   gpc1_1 gpc1_1_8332(
      {stage077[246]},
      {stage077[257]}
   );
   gpc1_1 gpc1_1_8333(
      {stage077[247]},
      {stage077[258]}
   );
   gpc1_1 gpc1_1_8334(
      {stage077[248]},
      {stage077[259]}
   );
   gpc1_1 gpc1_1_8335(
      {stage077[249]},
      {stage077[260]}
   );
   gpc1_1 gpc1_1_8336(
      {stage077[250]},
      {stage077[261]}
   );
   gpc1_1 gpc1_1_8337(
      {stage077[251]},
      {stage077[262]}
   );
   gpc1_1 gpc1_1_8338(
      {stage079[238]},
      {stage079[254]}
   );
   gpc1_1 gpc1_1_8339(
      {stage079[239]},
      {stage079[255]}
   );
   gpc1_1 gpc1_1_8340(
      {stage079[240]},
      {stage079[256]}
   );
   gpc1_1 gpc1_1_8341(
      {stage079[241]},
      {stage079[257]}
   );
   gpc606_5 gpc606_5_8342(
      {stage079[242], stage079[243], stage079[244], stage079[245], stage079[246], stage079[247]},
      {stage081[258], stage081[259], stage081[260], stage081[261], stage081[262], stage081[263]},
      {stage083[268], stage082[263], stage081[283], stage080[262], stage079[258]}
   );
   gpc615_5 gpc615_5_8343(
      {stage079[248], stage079[249], stage079[250], stage079[251], stage079[252]},
      {stage080[253]},
      {stage081[264], stage081[265], stage081[266], stage081[267], stage081[268], stage081[269]},
      {stage083[269], stage082[264], stage081[284], stage080[263], stage079[259]}
   );
   gpc1_1 gpc1_1_8344(
      {stage080[254]},
      {stage080[264]}
   );
   gpc606_5 gpc606_5_8345(
      {stage080[255], stage080[256], stage080[257], stage080[258], stage080[259], stage080[260]},
      {stage082[255], stage082[256], stage082[257], stage082[258], stage082[259], stage082[260]},
      {stage084[240], stage083[270], stage082[265], stage081[285], stage080[265]}
   );
   gpc1_1 gpc1_1_8346(
      {stage081[270]},
      {stage081[286]}
   );
   gpc1_1 gpc1_1_8347(
      {stage081[271]},
      {stage081[287]}
   );
   gpc1_1 gpc1_1_8348(
      {stage081[272]},
      {stage081[288]}
   );
   gpc1_1 gpc1_1_8349(
      {stage081[273]},
      {stage081[289]}
   );
   gpc1_1 gpc1_1_8350(
      {stage081[274]},
      {stage081[290]}
   );
   gpc1_1 gpc1_1_8351(
      {stage081[275]},
      {stage081[291]}
   );
   gpc207_4 gpc207_4_8352(
      {stage081[276], stage081[277], stage081[278], stage081[279], stage081[280], stage081[281], stage081[282]},
      {stage083[261], stage083[262]},
      {stage084[241], stage083[271], stage082[266], stage081[292]}
   );
   gpc1_1 gpc1_1_8353(
      {stage082[261]},
      {stage082[267]}
   );
   gpc1_1 gpc1_1_8354(
      {stage082[262]},
      {stage082[268]}
   );
   gpc1_1 gpc1_1_8355(
      {stage083[263]},
      {stage083[272]}
   );
   gpc1_1 gpc1_1_8356(
      {stage083[264]},
      {stage083[273]}
   );
   gpc1_1 gpc1_1_8357(
      {stage083[265]},
      {stage083[274]}
   );
   gpc1_1 gpc1_1_8358(
      {stage083[266]},
      {stage083[275]}
   );
   gpc1_1 gpc1_1_8359(
      {stage083[267]},
      {stage083[276]}
   );
   gpc606_5 gpc606_5_8360(
      {stage084[235], stage084[236], stage084[237], stage084[238], stage084[239], 1'h0},
      {stage086[271], stage086[272], stage086[273], stage086[274], stage086[275], stage086[276]},
      {stage088[274], stage087[237], stage086[284], stage085[274], stage084[242]}
   );
   gpc615_5 gpc615_5_8361(
      {stage085[265], stage085[266], stage085[267], stage085[268], stage085[269]},
      {stage086[277]},
      {stage087[223], stage087[224], stage087[225], stage087[226], stage087[227], stage087[228]},
      {stage089[266], stage088[275], stage087[238], stage086[285], stage085[275]}
   );
   gpc615_5 gpc615_5_8362(
      {stage085[270], stage085[271], stage085[272], stage085[273], 1'h0},
      {stage086[278]},
      {stage087[229], stage087[230], stage087[231], stage087[232], stage087[233], stage087[234]},
      {stage089[267], stage088[276], stage087[239], stage086[286], stage085[276]}
   );
   gpc1_1 gpc1_1_8363(
      {stage086[279]},
      {stage086[287]}
   );
   gpc1_1 gpc1_1_8364(
      {stage086[280]},
      {stage086[288]}
   );
   gpc1_1 gpc1_1_8365(
      {stage086[281]},
      {stage086[289]}
   );
   gpc1_1 gpc1_1_8366(
      {stage086[282]},
      {stage086[290]}
   );
   gpc1_1 gpc1_1_8367(
      {stage086[283]},
      {stage086[291]}
   );
   gpc1_1 gpc1_1_8368(
      {stage087[235]},
      {stage087[240]}
   );
   gpc1_1 gpc1_1_8369(
      {stage087[236]},
      {stage087[241]}
   );
   gpc1_1 gpc1_1_8370(
      {stage088[264]},
      {stage088[277]}
   );
   gpc1_1 gpc1_1_8371(
      {stage088[265]},
      {stage088[278]}
   );
   gpc1_1 gpc1_1_8372(
      {stage088[266]},
      {stage088[279]}
   );
   gpc1_1 gpc1_1_8373(
      {stage088[267]},
      {stage088[280]}
   );
   gpc606_5 gpc606_5_8374(
      {stage088[268], stage088[269], stage088[270], stage088[271], stage088[272], stage088[273]},
      {stage090[231], stage090[232], stage090[233], stage090[234], stage090[235], stage090[236]},
      {stage092[248], stage091[330], stage090[245], stage089[268], stage088[281]}
   );
   gpc1_1 gpc1_1_8375(
      {stage089[247]},
      {stage089[269]}
   );
   gpc606_5 gpc606_5_8376(
      {stage089[248], stage089[249], stage089[250], stage089[251], stage089[252], stage089[253]},
      {stage091[302], stage091[303], stage091[304], stage091[305], stage091[306], stage091[307]},
      {stage093[233], stage092[249], stage091[331], stage090[246], stage089[270]}
   );
   gpc606_5 gpc606_5_8377(
      {stage089[254], stage089[255], stage089[256], stage089[257], stage089[258], stage089[259]},
      {stage091[308], stage091[309], stage091[310], stage091[311], stage091[312], stage091[313]},
      {stage093[234], stage092[250], stage091[332], stage090[247], stage089[271]}
   );
   gpc606_5 gpc606_5_8378(
      {stage089[260], stage089[261], stage089[262], stage089[263], stage089[264], stage089[265]},
      {stage091[314], stage091[315], stage091[316], stage091[317], stage091[318], stage091[319]},
      {stage093[235], stage092[251], stage091[333], stage090[248], stage089[272]}
   );
   gpc1_1 gpc1_1_8379(
      {stage090[237]},
      {stage090[249]}
   );
   gpc1_1 gpc1_1_8380(
      {stage090[238]},
      {stage090[250]}
   );
   gpc1_1 gpc1_1_8381(
      {stage090[239]},
      {stage090[251]}
   );
   gpc615_5 gpc615_5_8382(
      {stage090[240], stage090[241], stage090[242], stage090[243], stage090[244]},
      {stage091[320]},
      {stage092[241], stage092[242], stage092[243], stage092[244], stage092[245], stage092[246]},
      {stage094[240], stage093[236], stage092[252], stage091[334], stage090[252]}
   );
   gpc1_1 gpc1_1_8383(
      {stage091[321]},
      {stage091[335]}
   );
   gpc1_1 gpc1_1_8384(
      {stage091[322]},
      {stage091[336]}
   );
   gpc1_1 gpc1_1_8385(
      {stage091[323]},
      {stage091[337]}
   );
   gpc606_5 gpc606_5_8386(
      {stage091[324], stage091[325], stage091[326], stage091[327], stage091[328], stage091[329]},
      {stage093[221], stage093[222], stage093[223], stage093[224], stage093[225], stage093[226]},
      {stage095[221], stage094[241], stage093[237], stage092[253], stage091[338]}
   );
   gpc1_1 gpc1_1_8387(
      {stage092[247]},
      {stage092[254]}
   );
   gpc606_5 gpc606_5_8388(
      {stage093[227], stage093[228], stage093[229], stage093[230], stage093[231], stage093[232]},
      {stage095[214], stage095[215], stage095[216], stage095[217], stage095[218], stage095[219]},
      {stage097[225], stage096[241], stage095[222], stage094[242], stage093[238]}
   );
   gpc606_5 gpc606_5_8389(
      {stage094[236], stage094[237], stage094[238], stage094[239], 1'h0, 1'h0},
      {stage096[231], stage096[232], stage096[233], stage096[234], stage096[235], stage096[236]},
      {stage098[239], stage097[226], stage096[242], stage095[223], stage094[243]}
   );
   gpc1_1 gpc1_1_8390(
      {stage095[220]},
      {stage095[224]}
   );
   gpc606_5 gpc606_5_8391(
      {stage096[237], stage096[238], stage096[239], stage096[240], 1'h0, 1'h0},
      {stage098[226], stage098[227], stage098[228], stage098[229], stage098[230], stage098[231]},
      {stage100[225], stage099[290], stage098[240], stage097[227], stage096[243]}
   );
   gpc615_5 gpc615_5_8392(
      {stage097[220], stage097[221], stage097[222], stage097[223], stage097[224]},
      {stage098[232]},
      {stage099[280], stage099[281], stage099[282], stage099[283], stage099[284], stage099[285]},
      {stage101[260], stage100[226], stage099[291], stage098[241], stage097[228]}
   );
   gpc1_1 gpc1_1_8393(
      {stage098[233]},
      {stage098[242]}
   );
   gpc615_5 gpc615_5_8394(
      {stage098[234], stage098[235], stage098[236], stage098[237], stage098[238]},
      {stage099[286]},
      {stage100[218], stage100[219], stage100[220], stage100[221], stage100[222], stage100[223]},
      {stage102[244], stage101[261], stage100[227], stage099[292], stage098[243]}
   );
   gpc1_1 gpc1_1_8395(
      {stage099[287]},
      {stage099[293]}
   );
   gpc1_1 gpc1_1_8396(
      {stage099[288]},
      {stage099[294]}
   );
   gpc1_1 gpc1_1_8397(
      {stage099[289]},
      {stage099[295]}
   );
   gpc1_1 gpc1_1_8398(
      {stage100[224]},
      {stage100[228]}
   );
   gpc1_1 gpc1_1_8399(
      {stage101[253]},
      {stage101[262]}
   );
   gpc1_1 gpc1_1_8400(
      {stage101[254]},
      {stage101[263]}
   );
   gpc615_5 gpc615_5_8401(
      {stage101[255], stage101[256], stage101[257], stage101[258], stage101[259]},
      {stage102[235]},
      {stage103[237], stage103[238], stage103[239], stage103[240], stage103[241], stage103[242]},
      {stage105[223], stage104[262], stage103[249], stage102[245], stage101[264]}
   );
   gpc1_1 gpc1_1_8402(
      {stage102[236]},
      {stage102[246]}
   );
   gpc1_1 gpc1_1_8403(
      {stage102[237]},
      {stage102[247]}
   );
   gpc1406_5 gpc1406_5_8404(
      {stage102[238], stage102[239], stage102[240], stage102[241], stage102[242], stage102[243]},
      {stage104[257], stage104[258], stage104[259], stage104[260]},
      {stage105[217]},
      {stage106[253], stage105[224], stage104[263], stage103[250], stage102[248]}
   );
   gpc1_1 gpc1_1_8405(
      {stage103[243]},
      {stage103[251]}
   );
   gpc1_1 gpc1_1_8406(
      {stage103[244]},
      {stage103[252]}
   );
   gpc1_1 gpc1_1_8407(
      {stage103[245]},
      {stage103[253]}
   );
   gpc623_5 gpc623_5_8408(
      {stage103[246], stage103[247], stage103[248]},
      {stage104[261], 1'h0},
      {stage105[218], stage105[219], stage105[220], stage105[221], stage105[222], 1'h0},
      {stage107[255], stage106[254], stage105[225], stage104[264], stage103[254]}
   );
   gpc615_5 gpc615_5_8409(
      {stage106[248], stage106[249], stage106[250], stage106[251], stage106[252]},
      {stage107[248]},
      {stage108[247], stage108[248], stage108[249], stage108[250], stage108[251], stage108[252]},
      {stage110[264], stage109[232], stage108[259], stage107[256], stage106[255]}
   );
   gpc1_1 gpc1_1_8410(
      {stage107[249]},
      {stage107[257]}
   );
   gpc1_1 gpc1_1_8411(
      {stage107[250]},
      {stage107[258]}
   );
   gpc1_1 gpc1_1_8412(
      {stage107[251]},
      {stage107[259]}
   );
   gpc1343_5 gpc1343_5_8413(
      {stage107[252], stage107[253], stage107[254]},
      {stage108[253], stage108[254], stage108[255], stage108[256]},
      {stage109[224], stage109[225], stage109[226]},
      {stage110[256]},
      {stage111[260], stage110[265], stage109[233], stage108[260], stage107[260]}
   );
   gpc1_1 gpc1_1_8414(
      {stage108[257]},
      {stage108[261]}
   );
   gpc1_1 gpc1_1_8415(
      {stage108[258]},
      {stage108[262]}
   );
   gpc615_5 gpc615_5_8416(
      {stage109[227], stage109[228], stage109[229], stage109[230], stage109[231]},
      {stage110[257]},
      {stage111[254], stage111[255], stage111[256], stage111[257], stage111[258], stage111[259]},
      {stage113[237], stage112[235], stage111[261], stage110[266], stage109[234]}
   );
   gpc606_5 gpc606_5_8417(
      {stage110[258], stage110[259], stage110[260], stage110[261], stage110[262], stage110[263]},
      {stage112[227], stage112[228], stage112[229], stage112[230], stage112[231], stage112[232]},
      {stage114[239], stage113[238], stage112[236], stage111[262], stage110[267]}
   );
   gpc1_1 gpc1_1_8418(
      {stage112[233]},
      {stage112[237]}
   );
   gpc1_1 gpc1_1_8419(
      {stage112[234]},
      {stage112[238]}
   );
   gpc1406_5 gpc1406_5_8420(
      {stage113[226], stage113[227], stage113[228], stage113[229], stage113[230], stage113[231]},
      {stage115[252], stage115[253], stage115[254], stage115[255]},
      {stage116[231]},
      {stage117[253], stage116[238], stage115[259], stage114[240], stage113[239]}
   );
   gpc1406_5 gpc1406_5_8421(
      {stage113[232], stage113[233], stage113[234], stage113[235], stage113[236], 1'h0},
      {stage115[256], stage115[257], stage115[258], 1'h0},
      {stage116[232]},
      {stage117[254], stage116[239], stage115[260], stage114[241], stage113[240]}
   );
   gpc1_1 gpc1_1_8422(
      {stage114[234]},
      {stage114[242]}
   );
   gpc1_1 gpc1_1_8423(
      {stage114[235]},
      {stage114[243]}
   );
   gpc1_1 gpc1_1_8424(
      {stage114[236]},
      {stage114[244]}
   );
   gpc1_1 gpc1_1_8425(
      {stage114[237]},
      {stage114[245]}
   );
   gpc1_1 gpc1_1_8426(
      {stage114[238]},
      {stage114[246]}
   );
   gpc2135_5 gpc2135_5_8427(
      {stage116[233], stage116[234], stage116[235], stage116[236], stage116[237]},
      {stage117[244], stage117[245], stage117[246]},
      {stage118[248]},
      {stage119[220], stage119[221]},
      {stage120[251], stage119[232], stage118[257], stage117[255], stage116[240]}
   );
   gpc615_5 gpc615_5_8428(
      {stage117[247], stage117[248], stage117[249], stage117[250], stage117[251]},
      {stage118[249]},
      {stage119[222], stage119[223], stage119[224], stage119[225], stage119[226], stage119[227]},
      {stage121[225], stage120[252], stage119[233], stage118[258], stage117[256]}
   );
   gpc1343_5 gpc1343_5_8429(
      {stage117[252], 1'h0, 1'h0},
      {stage118[250], stage118[251], stage118[252], stage118[253]},
      {stage119[228], stage119[229], stage119[230]},
      {stage120[245]},
      {stage121[226], stage120[253], stage119[234], stage118[259], stage117[257]}
   );
   gpc1_1 gpc1_1_8430(
      {stage118[254]},
      {stage118[260]}
   );
   gpc1_1 gpc1_1_8431(
      {stage118[255]},
      {stage118[261]}
   );
   gpc1_1 gpc1_1_8432(
      {stage118[256]},
      {stage118[262]}
   );
   gpc1_1 gpc1_1_8433(
      {stage119[231]},
      {stage119[235]}
   );
   gpc615_5 gpc615_5_8434(
      {stage120[246], stage120[247], stage120[248], stage120[249], stage120[250]},
      {stage121[217]},
      {stage122[235], stage122[236], stage122[237], stage122[238], stage122[239], stage122[240]},
      {stage124[229], stage123[318], stage122[243], stage121[227], stage120[254]}
   );
   gpc1_1 gpc1_1_8435(
      {stage121[218]},
      {stage121[228]}
   );
   gpc1_1 gpc1_1_8436(
      {stage121[219]},
      {stage121[229]}
   );
   gpc1_1 gpc1_1_8437(
      {stage121[220]},
      {stage121[230]}
   );
   gpc1_1 gpc1_1_8438(
      {stage121[221]},
      {stage121[231]}
   );
   gpc1_1 gpc1_1_8439(
      {stage121[222]},
      {stage121[232]}
   );
   gpc1_1 gpc1_1_8440(
      {stage121[223]},
      {stage121[233]}
   );
   gpc1_1 gpc1_1_8441(
      {stage121[224]},
      {stage121[234]}
   );
   gpc1_1 gpc1_1_8442(
      {stage122[241]},
      {stage122[244]}
   );
   gpc1_1 gpc1_1_8443(
      {stage122[242]},
      {stage122[245]}
   );
   gpc1_1 gpc1_1_8444(
      {stage123[306]},
      {stage123[319]}
   );
   gpc1_1 gpc1_1_8445(
      {stage123[307]},
      {stage123[320]}
   );
   gpc1_1 gpc1_1_8446(
      {stage123[308]},
      {stage123[321]}
   );
   gpc1_1 gpc1_1_8447(
      {stage123[309]},
      {stage123[322]}
   );
   gpc1_1 gpc1_1_8448(
      {stage123[310]},
      {stage123[323]}
   );
   gpc1_1 gpc1_1_8449(
      {stage123[311]},
      {stage123[324]}
   );
   gpc606_5 gpc606_5_8450(
      {stage123[312], stage123[313], stage123[314], stage123[315], stage123[316], stage123[317]},
      {stage125[263], stage125[264], stage125[265], stage125[266], stage125[267], stage125[268]},
      {stage127[281], stage126[277], stage125[280], stage124[230], stage123[325]}
   );
   gpc1_1 gpc1_1_8451(
      {stage124[224]},
      {stage124[231]}
   );
   gpc1_1 gpc1_1_8452(
      {stage124[225]},
      {stage124[232]}
   );
   gpc1_1 gpc1_1_8453(
      {stage124[226]},
      {stage124[233]}
   );
   gpc1_1 gpc1_1_8454(
      {stage124[227]},
      {stage124[234]}
   );
   gpc1_1 gpc1_1_8455(
      {stage124[228]},
      {stage124[235]}
   );
   gpc606_5 gpc606_5_8456(
      {stage125[269], stage125[270], stage125[271], stage125[272], stage125[273], stage125[274]},
      {stage127[268], stage127[269], stage127[270], stage127[271], stage127[272], stage127[273]},
      {stage129[66], stage128[83], stage127[282], stage126[278], stage125[281]}
   );
   gpc1325_5 gpc1325_5_8457(
      {stage125[275], stage125[276], stage125[277], stage125[278], stage125[279]},
      {stage126[263], stage126[264]},
      {stage127[274], stage127[275], stage127[276]},
      {stage128[72]},
      {stage129[67], stage128[84], stage127[283], stage126[279], stage125[282]}
   );
   gpc1_1 gpc1_1_8458(
      {stage126[265]},
      {stage126[280]}
   );
   gpc1_1 gpc1_1_8459(
      {stage126[266]},
      {stage126[281]}
   );
   gpc615_5 gpc615_5_8460(
      {stage126[267], stage126[268], stage126[269], stage126[270], stage126[271]},
      {stage127[277]},
      {stage128[73], stage128[74], stage128[75], stage128[76], stage128[77], stage128[78]},
      {stage130[14], stage129[68], stage128[85], stage127[284], stage126[282]}
   );
   gpc615_5 gpc615_5_8461(
      {stage126[272], stage126[273], stage126[274], stage126[275], stage126[276]},
      {stage127[278]},
      {stage128[79], stage128[80], stage128[81], stage128[82], 1'h0, 1'h0},
      {stage130[15], stage129[69], stage128[86], stage127[285], stage126[283]}
   );
   gpc1_1 gpc1_1_8462(
      {stage127[279]},
      {stage127[286]}
   );
   gpc1_1 gpc1_1_8463(
      {stage127[280]},
      {stage127[287]}
   );
   gpc1_1 gpc1_1_8464(
      {stage129[56]},
      {stage129[70]}
   );
   gpc1_1 gpc1_1_8465(
      {stage129[57]},
      {stage129[71]}
   );
   gpc1_1 gpc1_1_8466(
      {stage129[58]},
      {stage129[72]}
   );
   gpc1_1 gpc1_1_8467(
      {stage129[59]},
      {stage129[73]}
   );
   gpc1_1 gpc1_1_8468(
      {stage129[60]},
      {stage129[74]}
   );
   gpc1_1 gpc1_1_8469(
      {stage129[61]},
      {stage129[75]}
   );
   gpc1_1 gpc1_1_8470(
      {stage129[62]},
      {stage129[76]}
   );
   gpc1_1 gpc1_1_8471(
      {stage129[63]},
      {stage129[77]}
   );
   gpc1_1 gpc1_1_8472(
      {stage129[64]},
      {stage129[78]}
   );
   gpc1_1 gpc1_1_8473(
      {stage129[65]},
      {stage129[79]}
   );
   gpc207_4 gpc207_4_8474(
      {stage130[9], stage130[10], stage130[11], stage130[12], stage130[13], 1'h0, 1'h0},
      {stage132[1], stage132[2]},
      {stage133[1], stage132[4], stage131[7], stage130[16]}
   );
   gpc1_1 gpc1_1_8475(
      {stage131[4]},
      {stage131[8]}
   );
   gpc1_1 gpc1_1_8476(
      {stage131[5]},
      {stage131[9]}
   );
   gpc1_1 gpc1_1_8477(
      {stage131[6]},
      {stage131[10]}
   );
   gpc1_1 gpc1_1_8478(
      {stage132[3]},
      {stage132[5]}
   );
   gpc1_1 gpc1_1_8479(
      {stage133[0]},
      {stage133[2]}
   );
   gpc1_1 gpc1_1_8480(
      {stage000[188]},
      {stage000[190]}
   );
   gpc1_1 gpc1_1_8481(
      {stage000[189]},
      {stage000[191]}
   );
   gpc1_1 gpc1_1_8482(
      {stage001[226]},
      {stage001[228]}
   );
   gpc1_1 gpc1_1_8483(
      {stage001[227]},
      {stage001[229]}
   );
   gpc1_1 gpc1_1_8484(
      {stage002[242]},
      {stage002[244]}
   );
   gpc1_1 gpc1_1_8485(
      {stage002[243]},
      {stage002[245]}
   );
   gpc615_5 gpc615_5_8486(
      {stage003[214], stage003[215], stage003[216], stage003[217], 1'h0},
      {stage004[263]},
      {stage005[277], stage005[278], stage005[279], stage005[280], 1'h0, 1'h0},
      {stage007[257], stage006[258], stage005[281], stage004[270], stage003[218]}
   );
   gpc1_1 gpc1_1_8487(
      {stage004[264]},
      {stage004[271]}
   );
   gpc1_1 gpc1_1_8488(
      {stage004[265]},
      {stage004[272]}
   );
   gpc1_1 gpc1_1_8489(
      {stage004[266]},
      {stage004[273]}
   );
   gpc1_1 gpc1_1_8490(
      {stage004[267]},
      {stage004[274]}
   );
   gpc1_1 gpc1_1_8491(
      {stage004[268]},
      {stage004[275]}
   );
   gpc1_1 gpc1_1_8492(
      {stage004[269]},
      {stage004[276]}
   );
   gpc207_4 gpc207_4_8493(
      {stage006[251], stage006[252], stage006[253], stage006[254], stage006[255], stage006[256], stage006[257]},
      {stage008[236], stage008[237]},
      {stage009[239], stage008[245], stage007[258], stage006[259]}
   );
   gpc7_3 gpc7_3_8494(
      {stage007[250], stage007[251], stage007[252], stage007[253], stage007[254], stage007[255], stage007[256]},
      {stage009[240], stage008[246], stage007[259]}
   );
   gpc207_4 gpc207_4_8495(
      {stage008[238], stage008[239], stage008[240], stage008[241], stage008[242], stage008[243], stage008[244]},
      {stage010[291], stage010[292]},
      {stage011[261], stage010[299], stage009[241], stage008[247]}
   );
   gpc1_1 gpc1_1_8496(
      {stage009[237]},
      {stage009[242]}
   );
   gpc1_1 gpc1_1_8497(
      {stage009[238]},
      {stage009[243]}
   );
   gpc606_5 gpc606_5_8498(
      {stage010[293], stage010[294], stage010[295], stage010[296], stage010[297], stage010[298]},
      {stage012[319], stage012[320], stage012[321], stage012[322], stage012[323], stage012[324]},
      {stage014[304], stage013[268], stage012[325], stage011[262], stage010[300]}
   );
   gpc1_1 gpc1_1_8499(
      {stage011[254]},
      {stage011[263]}
   );
   gpc1_1 gpc1_1_8500(
      {stage011[255]},
      {stage011[264]}
   );
   gpc615_5 gpc615_5_8501(
      {stage011[256], stage011[257], stage011[258], stage011[259], stage011[260]},
      {1'h0},
      {stage013[253], stage013[254], stage013[255], stage013[256], stage013[257], stage013[258]},
      {stage015[260], stage014[305], stage013[269], stage012[326], stage011[265]}
   );
   gpc1_1 gpc1_1_8502(
      {stage013[259]},
      {stage013[270]}
   );
   gpc1_1 gpc1_1_8503(
      {stage013[260]},
      {stage013[271]}
   );
   gpc1_1 gpc1_1_8504(
      {stage013[261]},
      {stage013[272]}
   );
   gpc606_5 gpc606_5_8505(
      {stage013[262], stage013[263], stage013[264], stage013[265], stage013[266], stage013[267]},
      {stage015[253], stage015[254], stage015[255], stage015[256], stage015[257], stage015[258]},
      {stage017[281], stage016[291], stage015[261], stage014[306], stage013[273]}
   );
   gpc1_1 gpc1_1_8506(
      {stage014[298]},
      {stage014[307]}
   );
   gpc615_5 gpc615_5_8507(
      {stage014[299], stage014[300], stage014[301], stage014[302], stage014[303]},
      {stage015[259]},
      {stage016[285], stage016[286], stage016[287], stage016[288], stage016[289], stage016[290]},
      {stage018[254], stage017[282], stage016[292], stage015[262], stage014[308]}
   );
   gpc1_1 gpc1_1_8508(
      {stage017[278]},
      {stage017[283]}
   );
   gpc1_1 gpc1_1_8509(
      {stage017[279]},
      {stage017[284]}
   );
   gpc1_1 gpc1_1_8510(
      {stage017[280]},
      {stage017[285]}
   );
   gpc615_5 gpc615_5_8511(
      {stage018[249], stage018[250], stage018[251], stage018[252], stage018[253]},
      {stage019[258]},
      {stage020[229], stage020[230], stage020[231], stage020[232], stage020[233], stage020[234]},
      {stage022[231], stage021[295], stage020[235], stage019[269], stage018[255]}
   );
   gpc1_1 gpc1_1_8512(
      {stage019[259]},
      {stage019[270]}
   );
   gpc1_1 gpc1_1_8513(
      {stage019[260]},
      {stage019[271]}
   );
   gpc1_1 gpc1_1_8514(
      {stage019[261]},
      {stage019[272]}
   );
   gpc1_1 gpc1_1_8515(
      {stage019[262]},
      {stage019[273]}
   );
   gpc1_1 gpc1_1_8516(
      {stage019[263]},
      {stage019[274]}
   );
   gpc1_1 gpc1_1_8517(
      {stage019[264]},
      {stage019[275]}
   );
   gpc1_1 gpc1_1_8518(
      {stage019[265]},
      {stage019[276]}
   );
   gpc1_1 gpc1_1_8519(
      {stage019[266]},
      {stage019[277]}
   );
   gpc1_1 gpc1_1_8520(
      {stage019[267]},
      {stage019[278]}
   );
   gpc1_1 gpc1_1_8521(
      {stage019[268]},
      {stage019[279]}
   );
   gpc1_1 gpc1_1_8522(
      {stage021[285]},
      {stage021[296]}
   );
   gpc1_1 gpc1_1_8523(
      {stage021[286]},
      {stage021[297]}
   );
   gpc1_1 gpc1_1_8524(
      {stage021[287]},
      {stage021[298]}
   );
   gpc1_1 gpc1_1_8525(
      {stage021[288]},
      {stage021[299]}
   );
   gpc606_5 gpc606_5_8526(
      {stage021[289], stage021[290], stage021[291], stage021[292], stage021[293], stage021[294]},
      {stage023[309], stage023[310], stage023[311], stage023[312], stage023[313], stage023[314]},
      {stage025[296], stage024[259], stage023[317], stage022[232], stage021[300]}
   );
   gpc1_1 gpc1_1_8527(
      {stage022[225]},
      {stage022[233]}
   );
   gpc615_5 gpc615_5_8528(
      {stage022[226], stage022[227], stage022[228], stage022[229], stage022[230]},
      {stage023[315]},
      {stage024[254], stage024[255], stage024[256], stage024[257], stage024[258], 1'h0},
      {stage026[243], stage025[297], stage024[260], stage023[318], stage022[234]}
   );
   gpc1_1 gpc1_1_8529(
      {stage023[316]},
      {stage023[319]}
   );
   gpc1_1 gpc1_1_8530(
      {stage025[292]},
      {stage025[298]}
   );
   gpc1_1 gpc1_1_8531(
      {stage025[293]},
      {stage025[299]}
   );
   gpc1_1 gpc1_1_8532(
      {stage025[294]},
      {stage025[300]}
   );
   gpc1_1 gpc1_1_8533(
      {stage025[295]},
      {stage025[301]}
   );
   gpc1_1 gpc1_1_8534(
      {stage026[240]},
      {stage026[244]}
   );
   gpc1_1 gpc1_1_8535(
      {stage026[241]},
      {stage026[245]}
   );
   gpc1_1 gpc1_1_8536(
      {stage026[242]},
      {stage026[246]}
   );
   gpc7_3 gpc7_3_8537(
      {stage027[235], stage027[236], stage027[237], stage027[238], stage027[239], 1'h0, 1'h0},
      {stage029[288], stage028[265], stage027[240]}
   );
   gpc1_1 gpc1_1_8538(
      {stage028[254]},
      {stage028[266]}
   );
   gpc1_1 gpc1_1_8539(
      {stage028[255]},
      {stage028[267]}
   );
   gpc1_1 gpc1_1_8540(
      {stage028[256]},
      {stage028[268]}
   );
   gpc1_1 gpc1_1_8541(
      {stage028[257]},
      {stage028[269]}
   );
   gpc1_1 gpc1_1_8542(
      {stage028[258]},
      {stage028[270]}
   );
   gpc606_5 gpc606_5_8543(
      {stage028[259], stage028[260], stage028[261], stage028[262], stage028[263], stage028[264]},
      {stage030[240], stage030[241], stage030[242], stage030[243], stage030[244], stage030[245]},
      {stage032[304], stage031[255], stage030[247], stage029[289], stage028[271]}
   );
   gpc1_1 gpc1_1_8544(
      {stage029[285]},
      {stage029[290]}
   );
   gpc1_1 gpc1_1_8545(
      {stage029[286]},
      {stage029[291]}
   );
   gpc1_1 gpc1_1_8546(
      {stage029[287]},
      {stage029[292]}
   );
   gpc1_1 gpc1_1_8547(
      {stage030[246]},
      {stage030[248]}
   );
   gpc7_3 gpc7_3_8548(
      {stage031[250], stage031[251], stage031[252], stage031[253], stage031[254], 1'h0, 1'h0},
      {stage033[296], stage032[305], stage031[256]}
   );
   gpc207_4 gpc207_4_8549(
      {stage032[298], stage032[299], stage032[300], stage032[301], stage032[302], stage032[303], 1'h0},
      {stage034[299], stage034[300]},
      {stage035[265], stage034[309], stage033[297], stage032[306]}
   );
   gpc1_1 gpc1_1_8550(
      {stage033[291]},
      {stage033[298]}
   );
   gpc1_1 gpc1_1_8551(
      {stage033[292]},
      {stage033[299]}
   );
   gpc1_1 gpc1_1_8552(
      {stage033[293]},
      {stage033[300]}
   );
   gpc1_1 gpc1_1_8553(
      {stage033[294]},
      {stage033[301]}
   );
   gpc1_1 gpc1_1_8554(
      {stage033[295]},
      {stage033[302]}
   );
   gpc1_1 gpc1_1_8555(
      {stage034[301]},
      {stage034[310]}
   );
   gpc1_1 gpc1_1_8556(
      {stage034[302]},
      {stage034[311]}
   );
   gpc1_1 gpc1_1_8557(
      {stage034[303]},
      {stage034[312]}
   );
   gpc615_5 gpc615_5_8558(
      {stage034[304], stage034[305], stage034[306], stage034[307], stage034[308]},
      {stage035[260]},
      {stage036[225], stage036[226], stage036[227], stage036[228], stage036[229], stage036[230]},
      {stage038[257], stage037[279], stage036[231], stage035[266], stage034[313]}
   );
   gpc615_5 gpc615_5_8559(
      {stage035[261], stage035[262], stage035[263], stage035[264], 1'h0},
      {1'h0},
      {stage037[271], stage037[272], stage037[273], stage037[274], stage037[275], stage037[276]},
      {stage039[256], stage038[258], stage037[280], stage036[232], stage035[267]}
   );
   gpc623_5 gpc623_5_8560(
      {stage037[277], stage037[278], 1'h0},
      {stage038[250], stage038[251]},
      {stage039[250], stage039[251], stage039[252], stage039[253], stage039[254], stage039[255]},
      {stage041[278], stage040[307], stage039[257], stage038[259], stage037[281]}
   );
   gpc606_5 gpc606_5_8561(
      {stage038[252], stage038[253], stage038[254], stage038[255], stage038[256], 1'h0},
      {stage040[301], stage040[302], stage040[303], stage040[304], stage040[305], stage040[306]},
      {stage042[296], stage041[279], stage040[308], stage039[258], stage038[260]}
   );
   gpc1_1 gpc1_1_8562(
      {stage041[267]},
      {stage041[280]}
   );
   gpc1_1 gpc1_1_8563(
      {stage041[268]},
      {stage041[281]}
   );
   gpc1_1 gpc1_1_8564(
      {stage041[269]},
      {stage041[282]}
   );
   gpc1_1 gpc1_1_8565(
      {stage041[270]},
      {stage041[283]}
   );
   gpc207_4 gpc207_4_8566(
      {stage041[271], stage041[272], stage041[273], stage041[274], stage041[275], stage041[276], stage041[277]},
      {stage043[217], stage043[218]},
      {stage044[229], stage043[221], stage042[297], stage041[284]}
   );
   gpc1325_5 gpc1325_5_8567(
      {stage042[291], stage042[292], stage042[293], stage042[294], stage042[295]},
      {stage043[219], stage043[220]},
      {stage044[226], stage044[227], stage044[228]},
      {stage045[272]},
      {stage046[279], stage045[274], stage044[230], stage043[222], stage042[298]}
   );
   gpc1_1 gpc1_1_8568(
      {stage045[273]},
      {stage045[275]}
   );
   gpc207_4 gpc207_4_8569(
      {stage046[272], stage046[273], stage046[274], stage046[275], stage046[276], stage046[277], stage046[278]},
      {stage048[336], stage048[337]},
      {stage049[258], stage048[346], stage047[237], stage046[280]}
   );
   gpc1415_5 gpc1415_5_8570(
      {stage047[232], stage047[233], stage047[234], stage047[235], stage047[236]},
      {stage048[338]},
      {stage049[255], stage049[256], stage049[257], 1'h0},
      {stage050[278]},
      {stage051[254], stage050[283], stage049[259], stage048[347], stage047[238]}
   );
   gpc207_4 gpc207_4_8571(
      {stage048[339], stage048[340], stage048[341], stage048[342], stage048[343], stage048[344], stage048[345]},
      {stage050[279], stage050[280]},
      {stage051[255], stage050[284], stage049[260], stage048[348]}
   );
   gpc1_1 gpc1_1_8572(
      {stage050[281]},
      {stage050[285]}
   );
   gpc1_1 gpc1_1_8573(
      {stage050[282]},
      {stage050[286]}
   );
   gpc1_1 gpc1_1_8574(
      {stage051[249]},
      {stage051[256]}
   );
   gpc1_1 gpc1_1_8575(
      {stage051[250]},
      {stage051[257]}
   );
   gpc1_1 gpc1_1_8576(
      {stage051[251]},
      {stage051[258]}
   );
   gpc1_1 gpc1_1_8577(
      {stage051[252]},
      {stage051[259]}
   );
   gpc1_1 gpc1_1_8578(
      {stage051[253]},
      {stage051[260]}
   );
   gpc1_1 gpc1_1_8579(
      {stage052[274]},
      {stage052[278]}
   );
   gpc1_1 gpc1_1_8580(
      {stage052[275]},
      {stage052[279]}
   );
   gpc1_1 gpc1_1_8581(
      {stage052[276]},
      {stage052[280]}
   );
   gpc1_1 gpc1_1_8582(
      {stage052[277]},
      {stage052[281]}
   );
   gpc606_5 gpc606_5_8583(
      {stage053[249], stage053[250], stage053[251], stage053[252], stage053[253], stage053[254]},
      {stage055[284], stage055[285], stage055[286], stage055[287], stage055[288], stage055[289]},
      {stage057[259], stage056[292], stage055[295], stage054[262], stage053[255]}
   );
   gpc7_3 gpc7_3_8584(
      {stage054[255], stage054[256], stage054[257], stage054[258], stage054[259], stage054[260], stage054[261]},
      {stage056[293], stage055[296], stage054[263]}
   );
   gpc1_1 gpc1_1_8585(
      {stage055[290]},
      {stage055[297]}
   );
   gpc1_1 gpc1_1_8586(
      {stage055[291]},
      {stage055[298]}
   );
   gpc1_1 gpc1_1_8587(
      {stage055[292]},
      {stage055[299]}
   );
   gpc1_1 gpc1_1_8588(
      {stage055[293]},
      {stage055[300]}
   );
   gpc1_1 gpc1_1_8589(
      {stage055[294]},
      {stage055[301]}
   );
   gpc606_5 gpc606_5_8590(
      {stage056[286], stage056[287], stage056[288], stage056[289], stage056[290], stage056[291]},
      {stage058[232], stage058[233], stage058[234], stage058[235], stage058[236], 1'h0},
      {stage060[247], stage059[321], stage058[237], stage057[260], stage056[294]}
   );
   gpc207_4 gpc207_4_8591(
      {stage057[252], stage057[253], stage057[254], stage057[255], stage057[256], stage057[257], stage057[258]},
      {stage059[313], stage059[314]},
      {stage060[248], stage059[322], stage058[238], stage057[261]}
   );
   gpc606_5 gpc606_5_8592(
      {stage059[315], stage059[316], stage059[317], stage059[318], stage059[319], stage059[320]},
      {stage061[276], stage061[277], stage061[278], stage061[279], stage061[280], 1'h0},
      {stage063[219], stage062[259], stage061[281], stage060[249], stage059[323]}
   );
   gpc1_1 gpc1_1_8593(
      {stage060[240]},
      {stage060[250]}
   );
   gpc606_5 gpc606_5_8594(
      {stage060[241], stage060[242], stage060[243], stage060[244], stage060[245], stage060[246]},
      {stage062[253], stage062[254], stage062[255], stage062[256], stage062[257], stage062[258]},
      {stage064[269], stage063[220], stage062[260], stage061[282], stage060[251]}
   );
   gpc1_1 gpc1_1_8595(
      {stage063[215]},
      {stage063[221]}
   );
   gpc1_1 gpc1_1_8596(
      {stage063[216]},
      {stage063[222]}
   );
   gpc1_1 gpc1_1_8597(
      {stage063[217]},
      {stage063[223]}
   );
   gpc1_1 gpc1_1_8598(
      {stage063[218]},
      {stage063[224]}
   );
   gpc606_5 gpc606_5_8599(
      {stage064[264], stage064[265], stage064[266], stage064[267], stage064[268], 1'h0},
      {stage066[286], stage066[287], stage066[288], stage066[289], 1'h0, 1'h0},
      {stage068[281], stage067[268], stage066[290], stage065[264], stage064[270]}
   );
   gpc1_1 gpc1_1_8600(
      {stage065[261]},
      {stage065[265]}
   );
   gpc1_1 gpc1_1_8601(
      {stage065[262]},
      {stage065[266]}
   );
   gpc1_1 gpc1_1_8602(
      {stage065[263]},
      {stage065[267]}
   );
   gpc606_5 gpc606_5_8603(
      {stage067[262], stage067[263], stage067[264], stage067[265], stage067[266], stage067[267]},
      {stage069[263], stage069[264], stage069[265], stage069[266], stage069[267], stage069[268]},
      {stage071[266], stage070[265], stage069[272], stage068[282], stage067[269]}
   );
   gpc1_1 gpc1_1_8604(
      {stage068[277]},
      {stage068[283]}
   );
   gpc1_1 gpc1_1_8605(
      {stage068[278]},
      {stage068[284]}
   );
   gpc1_1 gpc1_1_8606(
      {stage068[279]},
      {stage068[285]}
   );
   gpc1_1 gpc1_1_8607(
      {stage068[280]},
      {stage068[286]}
   );
   gpc1_1 gpc1_1_8608(
      {stage069[269]},
      {stage069[273]}
   );
   gpc1_1 gpc1_1_8609(
      {stage069[270]},
      {stage069[274]}
   );
   gpc1_1 gpc1_1_8610(
      {stage069[271]},
      {stage069[275]}
   );
   gpc1_1 gpc1_1_8611(
      {stage070[259]},
      {stage070[266]}
   );
   gpc1415_5 gpc1415_5_8612(
      {stage070[260], stage070[261], stage070[262], stage070[263], stage070[264]},
      {stage071[263]},
      {stage072[311], stage072[312], stage072[313], stage072[314]},
      {stage073[243]},
      {stage074[262], stage073[247], stage072[315], stage071[267], stage070[267]}
   );
   gpc1_1 gpc1_1_8613(
      {stage071[264]},
      {stage071[268]}
   );
   gpc1_1 gpc1_1_8614(
      {stage071[265]},
      {stage071[269]}
   );
   gpc1_1 gpc1_1_8615(
      {stage073[244]},
      {stage073[248]}
   );
   gpc1_1 gpc1_1_8616(
      {stage073[245]},
      {stage073[249]}
   );
   gpc1_1 gpc1_1_8617(
      {stage073[246]},
      {stage073[250]}
   );
   gpc1_1 gpc1_1_8618(
      {stage074[254]},
      {stage074[263]}
   );
   gpc1_1 gpc1_1_8619(
      {stage074[255]},
      {stage074[264]}
   );
   gpc1406_5 gpc1406_5_8620(
      {stage074[256], stage074[257], stage074[258], stage074[259], stage074[260], stage074[261]},
      {stage076[215], stage076[216], stage076[217], 1'h0},
      {stage077[252]},
      {stage078[235], stage077[263], stage076[218], stage075[212], stage074[265]}
   );
   gpc606_5 gpc606_5_8621(
      {stage075[209], stage075[210], stage075[211], 1'h0, 1'h0, 1'h0},
      {stage077[253], stage077[254], stage077[255], stage077[256], stage077[257], stage077[258]},
      {stage079[260], stage078[236], stage077[264], stage076[219], stage075[213]}
   );
   gpc1_1 gpc1_1_8622(
      {stage077[259]},
      {stage077[265]}
   );
   gpc1_1 gpc1_1_8623(
      {stage077[260]},
      {stage077[266]}
   );
   gpc1_1 gpc1_1_8624(
      {stage077[261]},
      {stage077[267]}
   );
   gpc1_1 gpc1_1_8625(
      {stage077[262]},
      {stage077[268]}
   );
   gpc1_1 gpc1_1_8626(
      {stage078[234]},
      {stage078[237]}
   );
   gpc1_1 gpc1_1_8627(
      {stage079[253]},
      {stage079[261]}
   );
   gpc606_5 gpc606_5_8628(
      {stage079[254], stage079[255], stage079[256], stage079[257], stage079[258], stage079[259]},
      {stage081[283], stage081[284], stage081[285], stage081[286], stage081[287], stage081[288]},
      {stage083[277], stage082[269], stage081[293], stage080[266], stage079[262]}
   );
   gpc615_5 gpc615_5_8629(
      {stage080[261], stage080[262], stage080[263], stage080[264], stage080[265]},
      {stage081[289]},
      {stage082[263], stage082[264], stage082[265], stage082[266], stage082[267], stage082[268]},
      {stage084[243], stage083[278], stage082[270], stage081[294], stage080[267]}
   );
   gpc1_1 gpc1_1_8630(
      {stage081[290]},
      {stage081[295]}
   );
   gpc1_1 gpc1_1_8631(
      {stage081[291]},
      {stage081[296]}
   );
   gpc1_1 gpc1_1_8632(
      {stage081[292]},
      {stage081[297]}
   );
   gpc1_1 gpc1_1_8633(
      {stage083[268]},
      {stage083[279]}
   );
   gpc1_1 gpc1_1_8634(
      {stage083[269]},
      {stage083[280]}
   );
   gpc207_4 gpc207_4_8635(
      {stage083[270], stage083[271], stage083[272], stage083[273], stage083[274], stage083[275], stage083[276]},
      {stage085[274], stage085[275]},
      {stage086[292], stage085[277], stage084[244], stage083[281]}
   );
   gpc1_1 gpc1_1_8636(
      {stage084[240]},
      {stage084[245]}
   );
   gpc1_1 gpc1_1_8637(
      {stage084[241]},
      {stage084[246]}
   );
   gpc1_1 gpc1_1_8638(
      {stage084[242]},
      {stage084[247]}
   );
   gpc1_1 gpc1_1_8639(
      {stage085[276]},
      {stage085[278]}
   );
   gpc1_1 gpc1_1_8640(
      {stage086[284]},
      {stage086[293]}
   );
   gpc1_1 gpc1_1_8641(
      {stage086[285]},
      {stage086[294]}
   );
   gpc606_5 gpc606_5_8642(
      {stage086[286], stage086[287], stage086[288], stage086[289], stage086[290], stage086[291]},
      {stage088[274], stage088[275], stage088[276], stage088[277], stage088[278], stage088[279]},
      {stage090[253], stage089[273], stage088[282], stage087[242], stage086[295]}
   );
   gpc606_5 gpc606_5_8643(
      {stage087[237], stage087[238], stage087[239], stage087[240], stage087[241], 1'h0},
      {stage089[266], stage089[267], stage089[268], stage089[269], stage089[270], stage089[271]},
      {stage091[339], stage090[254], stage089[274], stage088[283], stage087[243]}
   );
   gpc1_1 gpc1_1_8644(
      {stage088[280]},
      {stage088[284]}
   );
   gpc1_1 gpc1_1_8645(
      {stage088[281]},
      {stage088[285]}
   );
   gpc1_1 gpc1_1_8646(
      {stage089[272]},
      {stage089[275]}
   );
   gpc1_1 gpc1_1_8647(
      {stage090[245]},
      {stage090[255]}
   );
   gpc1_1 gpc1_1_8648(
      {stage090[246]},
      {stage090[256]}
   );
   gpc1_1 gpc1_1_8649(
      {stage090[247]},
      {stage090[257]}
   );
   gpc615_5 gpc615_5_8650(
      {stage090[248], stage090[249], stage090[250], stage090[251], stage090[252]},
      {stage091[330]},
      {stage092[248], stage092[249], stage092[250], stage092[251], stage092[252], stage092[253]},
      {stage094[244], stage093[239], stage092[255], stage091[340], stage090[258]}
   );
   gpc1_1 gpc1_1_8651(
      {stage091[331]},
      {stage091[341]}
   );
   gpc1_1 gpc1_1_8652(
      {stage091[332]},
      {stage091[342]}
   );
   gpc606_5 gpc606_5_8653(
      {stage091[333], stage091[334], stage091[335], stage091[336], stage091[337], stage091[338]},
      {stage093[233], stage093[234], stage093[235], stage093[236], stage093[237], stage093[238]},
      {stage095[225], stage094[245], stage093[240], stage092[256], stage091[343]}
   );
   gpc1_1 gpc1_1_8654(
      {stage092[254]},
      {stage092[257]}
   );
   gpc1_1 gpc1_1_8655(
      {stage094[240]},
      {stage094[246]}
   );
   gpc1_1 gpc1_1_8656(
      {stage094[241]},
      {stage094[247]}
   );
   gpc1_1 gpc1_1_8657(
      {stage094[242]},
      {stage094[248]}
   );
   gpc1_1 gpc1_1_8658(
      {stage094[243]},
      {stage094[249]}
   );
   gpc1_1 gpc1_1_8659(
      {stage095[221]},
      {stage095[226]}
   );
   gpc1_1 gpc1_1_8660(
      {stage095[222]},
      {stage095[227]}
   );
   gpc1_1 gpc1_1_8661(
      {stage095[223]},
      {stage095[228]}
   );
   gpc1_1 gpc1_1_8662(
      {stage095[224]},
      {stage095[229]}
   );
   gpc1_1 gpc1_1_8663(
      {stage096[241]},
      {stage096[244]}
   );
   gpc1_1 gpc1_1_8664(
      {stage096[242]},
      {stage096[245]}
   );
   gpc1_1 gpc1_1_8665(
      {stage096[243]},
      {stage096[246]}
   );
   gpc1_1 gpc1_1_8666(
      {stage097[225]},
      {stage097[229]}
   );
   gpc1_1 gpc1_1_8667(
      {stage097[226]},
      {stage097[230]}
   );
   gpc1_1 gpc1_1_8668(
      {stage097[227]},
      {stage097[231]}
   );
   gpc1_1 gpc1_1_8669(
      {stage097[228]},
      {stage097[232]}
   );
   gpc606_5 gpc606_5_8670(
      {stage098[239], stage098[240], stage098[241], stage098[242], stage098[243], 1'h0},
      {stage100[225], stage100[226], stage100[227], stage100[228], 1'h0, 1'h0},
      {stage102[249], stage101[265], stage100[229], stage099[296], stage098[244]}
   );
   gpc1_1 gpc1_1_8671(
      {stage099[290]},
      {stage099[297]}
   );
   gpc1_1 gpc1_1_8672(
      {stage099[291]},
      {stage099[298]}
   );
   gpc1_1 gpc1_1_8673(
      {stage099[292]},
      {stage099[299]}
   );
   gpc1_1 gpc1_1_8674(
      {stage099[293]},
      {stage099[300]}
   );
   gpc1_1 gpc1_1_8675(
      {stage099[294]},
      {stage099[301]}
   );
   gpc1_1 gpc1_1_8676(
      {stage099[295]},
      {stage099[302]}
   );
   gpc1_1 gpc1_1_8677(
      {stage101[260]},
      {stage101[266]}
   );
   gpc1_1 gpc1_1_8678(
      {stage101[261]},
      {stage101[267]}
   );
   gpc1_1 gpc1_1_8679(
      {stage101[262]},
      {stage101[268]}
   );
   gpc1_1 gpc1_1_8680(
      {stage101[263]},
      {stage101[269]}
   );
   gpc1_1 gpc1_1_8681(
      {stage101[264]},
      {stage101[270]}
   );
   gpc615_5 gpc615_5_8682(
      {stage102[244], stage102[245], stage102[246], stage102[247], stage102[248]},
      {stage103[249]},
      {stage104[262], stage104[263], stage104[264], 1'h0, 1'h0, 1'h0},
      {stage106[256], stage105[226], stage104[265], stage103[255], stage102[250]}
   );
   gpc1_1 gpc1_1_8683(
      {stage103[250]},
      {stage103[256]}
   );
   gpc1_1 gpc1_1_8684(
      {stage103[251]},
      {stage103[257]}
   );
   gpc1_1 gpc1_1_8685(
      {stage103[252]},
      {stage103[258]}
   );
   gpc1_1 gpc1_1_8686(
      {stage103[253]},
      {stage103[259]}
   );
   gpc1_1 gpc1_1_8687(
      {stage103[254]},
      {stage103[260]}
   );
   gpc1_1 gpc1_1_8688(
      {stage105[223]},
      {stage105[227]}
   );
   gpc1_1 gpc1_1_8689(
      {stage105[224]},
      {stage105[228]}
   );
   gpc1_1 gpc1_1_8690(
      {stage105[225]},
      {stage105[229]}
   );
   gpc1_1 gpc1_1_8691(
      {stage106[253]},
      {stage106[257]}
   );
   gpc1_1 gpc1_1_8692(
      {stage106[254]},
      {stage106[258]}
   );
   gpc1_1 gpc1_1_8693(
      {stage106[255]},
      {stage106[259]}
   );
   gpc1_1 gpc1_1_8694(
      {stage107[255]},
      {stage107[261]}
   );
   gpc1_1 gpc1_1_8695(
      {stage107[256]},
      {stage107[262]}
   );
   gpc1_1 gpc1_1_8696(
      {stage107[257]},
      {stage107[263]}
   );
   gpc1_1 gpc1_1_8697(
      {stage107[258]},
      {stage107[264]}
   );
   gpc1_1 gpc1_1_8698(
      {stage107[259]},
      {stage107[265]}
   );
   gpc1_1 gpc1_1_8699(
      {stage107[260]},
      {stage107[266]}
   );
   gpc2135_5 gpc2135_5_8700(
      {stage108[259], stage108[260], stage108[261], stage108[262], 1'h0},
      {stage109[232], stage109[233], stage109[234]},
      {stage110[264]},
      {stage111[260], stage111[261]},
      {stage112[239], stage111[263], stage110[268], stage109[235], stage108[263]}
   );
   gpc1_1 gpc1_1_8701(
      {stage110[265]},
      {stage110[269]}
   );
   gpc1_1 gpc1_1_8702(
      {stage110[266]},
      {stage110[270]}
   );
   gpc1_1 gpc1_1_8703(
      {stage110[267]},
      {stage110[271]}
   );
   gpc1_1 gpc1_1_8704(
      {stage111[262]},
      {stage111[264]}
   );
   gpc1_1 gpc1_1_8705(
      {stage112[235]},
      {stage112[240]}
   );
   gpc1_1 gpc1_1_8706(
      {stage112[236]},
      {stage112[241]}
   );
   gpc1_1 gpc1_1_8707(
      {stage112[237]},
      {stage112[242]}
   );
   gpc1_1 gpc1_1_8708(
      {stage112[238]},
      {stage112[243]}
   );
   gpc2135_5 gpc2135_5_8709(
      {stage113[237], stage113[238], stage113[239], stage113[240], 1'h0},
      {stage114[239], stage114[240], stage114[241]},
      {stage115[259]},
      {stage116[238], stage116[239]},
      {stage117[258], stage116[241], stage115[261], stage114[247], stage113[241]}
   );
   gpc1_1 gpc1_1_8710(
      {stage114[242]},
      {stage114[248]}
   );
   gpc1_1 gpc1_1_8711(
      {stage114[243]},
      {stage114[249]}
   );
   gpc1_1 gpc1_1_8712(
      {stage114[244]},
      {stage114[250]}
   );
   gpc1_1 gpc1_1_8713(
      {stage114[245]},
      {stage114[251]}
   );
   gpc1_1 gpc1_1_8714(
      {stage114[246]},
      {stage114[252]}
   );
   gpc1_1 gpc1_1_8715(
      {stage115[260]},
      {stage115[262]}
   );
   gpc1_1 gpc1_1_8716(
      {stage116[240]},
      {stage116[242]}
   );
   gpc1_1 gpc1_1_8717(
      {stage117[253]},
      {stage117[259]}
   );
   gpc1_1 gpc1_1_8718(
      {stage117[254]},
      {stage117[260]}
   );
   gpc1_1 gpc1_1_8719(
      {stage117[255]},
      {stage117[261]}
   );
   gpc1_1 gpc1_1_8720(
      {stage117[256]},
      {stage117[262]}
   );
   gpc1_1 gpc1_1_8721(
      {stage117[257]},
      {stage117[263]}
   );
   gpc606_5 gpc606_5_8722(
      {stage118[257], stage118[258], stage118[259], stage118[260], stage118[261], stage118[262]},
      {stage120[251], stage120[252], stage120[253], stage120[254], 1'h0, 1'h0},
      {stage122[246], stage121[235], stage120[255], stage119[236], stage118[263]}
   );
   gpc1_1 gpc1_1_8723(
      {stage119[232]},
      {stage119[237]}
   );
   gpc1_1 gpc1_1_8724(
      {stage119[233]},
      {stage119[238]}
   );
   gpc1_1 gpc1_1_8725(
      {stage119[234]},
      {stage119[239]}
   );
   gpc1_1 gpc1_1_8726(
      {stage119[235]},
      {stage119[240]}
   );
   gpc1_1 gpc1_1_8727(
      {stage121[225]},
      {stage121[236]}
   );
   gpc1_1 gpc1_1_8728(
      {stage121[226]},
      {stage121[237]}
   );
   gpc1_1 gpc1_1_8729(
      {stage121[227]},
      {stage121[238]}
   );
   gpc1_1 gpc1_1_8730(
      {stage121[228]},
      {stage121[239]}
   );
   gpc606_5 gpc606_5_8731(
      {stage121[229], stage121[230], stage121[231], stage121[232], stage121[233], stage121[234]},
      {stage123[318], stage123[319], stage123[320], stage123[321], stage123[322], stage123[323]},
      {stage125[283], stage124[236], stage123[326], stage122[247], stage121[240]}
   );
   gpc1325_5 gpc1325_5_8732(
      {stage122[243], stage122[244], stage122[245], 1'h0, 1'h0},
      {stage123[324], stage123[325]},
      {stage124[229], stage124[230], stage124[231]},
      {stage125[280]},
      {stage126[284], stage125[284], stage124[237], stage123[327], stage122[248]}
   );
   gpc2135_5 gpc2135_5_8733(
      {stage124[232], stage124[233], stage124[234], stage124[235], 1'h0},
      {stage125[281], stage125[282], 1'h0},
      {stage126[277]},
      {stage127[281], stage127[282]},
      {stage128[87], stage127[288], stage126[285], stage125[285], stage124[238]}
   );
   gpc606_5 gpc606_5_8734(
      {stage126[278], stage126[279], stage126[280], stage126[281], stage126[282], stage126[283]},
      {stage128[83], stage128[84], stage128[85], stage128[86], 1'h0, 1'h0},
      {stage130[17], stage129[80], stage128[88], stage127[289], stage126[286]}
   );
   gpc606_5 gpc606_5_8735(
      {stage127[283], stage127[284], stage127[285], stage127[286], stage127[287], 1'h0},
      {stage129[66], stage129[67], stage129[68], stage129[69], stage129[70], stage129[71]},
      {stage131[11], stage130[18], stage129[81], stage128[89], stage127[290]}
   );
   gpc1_1 gpc1_1_8736(
      {stage129[72]},
      {stage129[82]}
   );
   gpc1_1 gpc1_1_8737(
      {stage129[73]},
      {stage129[83]}
   );
   gpc1_1 gpc1_1_8738(
      {stage129[74]},
      {stage129[84]}
   );
   gpc2135_5 gpc2135_5_8739(
      {stage129[75], stage129[76], stage129[77], stage129[78], stage129[79]},
      {stage130[14], stage130[15], stage130[16]},
      {stage131[7]},
      {stage132[4], stage132[5]},
      {stage133[3], stage132[6], stage131[12], stage130[19], stage129[85]}
   );
   gpc1_1 gpc1_1_8740(
      {stage131[8]},
      {stage131[13]}
   );
   gpc1_1 gpc1_1_8741(
      {stage131[9]},
      {stage131[14]}
   );
   gpc1_1 gpc1_1_8742(
      {stage131[10]},
      {stage131[15]}
   );
   gpc1_1 gpc1_1_8743(
      {stage133[1]},
      {stage133[4]}
   );
   gpc1_1 gpc1_1_8744(
      {stage133[2]},
      {stage133[5]}
   );
   gpc1_1 gpc1_1_8745(
      {stage000[190]},
      {stage000[192]}
   );
   gpc1_1 gpc1_1_8746(
      {stage000[191]},
      {stage000[193]}
   );
   gpc1_1 gpc1_1_8747(
      {stage001[228]},
      {stage001[230]}
   );
   gpc1_1 gpc1_1_8748(
      {stage001[229]},
      {stage001[231]}
   );
   gpc1_1 gpc1_1_8749(
      {stage002[244]},
      {stage002[246]}
   );
   gpc1_1 gpc1_1_8750(
      {stage002[245]},
      {stage002[247]}
   );
   gpc1_1 gpc1_1_8751(
      {stage003[218]},
      {stage003[219]}
   );
   gpc207_4 gpc207_4_8752(
      {stage004[270], stage004[271], stage004[272], stage004[273], stage004[274], stage004[275], stage004[276]},
      {stage006[258], stage006[259]},
      {stage007[260], stage006[260], stage005[282], stage004[277]}
   );
   gpc1_1 gpc1_1_8753(
      {stage005[281]},
      {stage005[283]}
   );
   gpc23_3 gpc23_3_8754(
      {stage007[257], stage007[258], stage007[259]},
      {stage008[245], stage008[246]},
      {stage009[244], stage008[248], stage007[261]}
   );
   gpc1_1 gpc1_1_8755(
      {stage008[247]},
      {stage008[249]}
   );
   gpc215_4 gpc215_4_8756(
      {stage009[239], stage009[240], stage009[241], stage009[242], stage009[243]},
      {stage010[299]},
      {stage011[261], stage011[262]},
      {stage012[327], stage011[266], stage010[301], stage009[245]}
   );
   gpc1_1 gpc1_1_8757(
      {stage010[300]},
      {stage010[302]}
   );
   gpc623_5 gpc623_5_8758(
      {stage011[263], stage011[264], stage011[265]},
      {stage012[325], stage012[326]},
      {stage013[268], stage013[269], stage013[270], stage013[271], stage013[272], stage013[273]},
      {stage015[263], stage014[309], stage013[274], stage012[328], stage011[267]}
   );
   gpc135_4 gpc135_4_8759(
      {stage014[304], stage014[305], stage014[306], stage014[307], stage014[308]},
      {stage015[260], stage015[261], stage015[262]},
      {stage016[291]},
      {stage017[286], stage016[293], stage015[264], stage014[310]}
   );
   gpc1_1 gpc1_1_8760(
      {stage016[292]},
      {stage016[294]}
   );
   gpc615_5 gpc615_5_8761(
      {stage017[281], stage017[282], stage017[283], stage017[284], stage017[285]},
      {stage018[254]},
      {stage019[269], stage019[270], stage019[271], stage019[272], stage019[273], stage019[274]},
      {stage021[301], stage020[236], stage019[280], stage018[256], stage017[287]}
   );
   gpc1_1 gpc1_1_8762(
      {stage018[255]},
      {stage018[257]}
   );
   gpc615_5 gpc615_5_8763(
      {stage019[275], stage019[276], stage019[277], stage019[278], stage019[279]},
      {stage020[235]},
      {stage021[295], stage021[296], stage021[297], stage021[298], stage021[299], stage021[300]},
      {stage023[320], stage022[235], stage021[302], stage020[237], stage019[281]}
   );
   gpc135_4 gpc135_4_8764(
      {stage022[231], stage022[232], stage022[233], stage022[234], 1'h0},
      {stage023[317], stage023[318], stage023[319]},
      {stage024[259]},
      {stage025[302], stage024[261], stage023[321], stage022[236]}
   );
   gpc1_1 gpc1_1_8765(
      {stage024[260]},
      {stage024[262]}
   );
   gpc7_3 gpc7_3_8766(
      {stage025[296], stage025[297], stage025[298], stage025[299], stage025[300], stage025[301], 1'h0},
      {stage027[241], stage026[247], stage025[303]}
   );
   gpc615_5 gpc615_5_8767(
      {stage026[243], stage026[244], stage026[245], stage026[246], 1'h0},
      {stage027[240]},
      {stage028[265], stage028[266], stage028[267], stage028[268], stage028[269], stage028[270]},
      {stage030[249], stage029[293], stage028[272], stage027[242], stage026[248]}
   );
   gpc1_1 gpc1_1_8768(
      {stage028[271]},
      {stage028[273]}
   );
   gpc2135_5 gpc2135_5_8769(
      {stage029[288], stage029[289], stage029[290], stage029[291], stage029[292]},
      {stage030[247], stage030[248], 1'h0},
      {stage031[255]},
      {stage032[304], stage032[305]},
      {stage033[303], stage032[307], stage031[257], stage030[250], stage029[294]}
   );
   gpc1_1 gpc1_1_8770(
      {stage031[256]},
      {stage031[258]}
   );
   gpc1_1 gpc1_1_8771(
      {stage032[306]},
      {stage032[308]}
   );
   gpc7_3 gpc7_3_8772(
      {stage033[296], stage033[297], stage033[298], stage033[299], stage033[300], stage033[301], stage033[302]},
      {stage035[268], stage034[314], stage033[304]}
   );
   gpc135_4 gpc135_4_8773(
      {stage034[309], stage034[310], stage034[311], stage034[312], stage034[313]},
      {stage035[265], stage035[266], stage035[267]},
      {stage036[231]},
      {stage037[282], stage036[233], stage035[269], stage034[315]}
   );
   gpc1_1 gpc1_1_8774(
      {stage036[232]},
      {stage036[234]}
   );
   gpc1343_5 gpc1343_5_8775(
      {stage037[279], stage037[280], stage037[281]},
      {stage038[257], stage038[258], stage038[259], stage038[260]},
      {stage039[256], stage039[257], stage039[258]},
      {stage040[307]},
      {stage041[285], stage040[309], stage039[259], stage038[261], stage037[283]}
   );
   gpc1_1 gpc1_1_8776(
      {stage040[308]},
      {stage040[310]}
   );
   gpc207_4 gpc207_4_8777(
      {stage041[278], stage041[279], stage041[280], stage041[281], stage041[282], stage041[283], stage041[284]},
      {stage043[221], stage043[222]},
      {stage044[231], stage043[223], stage042[299], stage041[286]}
   );
   gpc615_5 gpc615_5_8778(
      {stage042[296], stage042[297], stage042[298], 1'h0, 1'h0},
      {1'h0},
      {stage044[229], stage044[230], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage046[281], stage045[276], stage044[232], stage043[224], stage042[300]}
   );
   gpc2135_5 gpc2135_5_8779(
      {stage045[274], stage045[275], 1'h0, 1'h0, 1'h0},
      {stage046[279], stage046[280], 1'h0},
      {stage047[237]},
      {stage048[346], stage048[347]},
      {stage049[261], stage048[349], stage047[239], stage046[282], stage045[277]}
   );
   gpc1_1 gpc1_1_8780(
      {stage047[238]},
      {stage047[240]}
   );
   gpc1_1 gpc1_1_8781(
      {stage048[348]},
      {stage048[350]}
   );
   gpc623_5 gpc623_5_8782(
      {stage049[258], stage049[259], stage049[260]},
      {stage050[283], stage050[284]},
      {stage051[254], stage051[255], stage051[256], stage051[257], stage051[258], stage051[259]},
      {stage053[256], stage052[282], stage051[261], stage050[287], stage049[262]}
   );
   gpc1415_5 gpc1415_5_8783(
      {stage050[285], stage050[286], 1'h0, 1'h0, 1'h0},
      {stage051[260]},
      {stage052[278], stage052[279], stage052[280], stage052[281]},
      {stage053[255]},
      {stage054[264], stage053[257], stage052[283], stage051[262], stage050[288]}
   );
   gpc223_4 gpc223_4_8784(
      {stage054[262], stage054[263], 1'h0},
      {stage055[295], stage055[296]},
      {stage056[292], stage056[293]},
      {stage057[262], stage056[295], stage055[302], stage054[265]}
   );
   gpc1325_5 gpc1325_5_8785(
      {stage055[297], stage055[298], stage055[299], stage055[300], stage055[301]},
      {stage056[294], 1'h0},
      {stage057[259], stage057[260], stage057[261]},
      {stage058[237]},
      {stage059[324], stage058[239], stage057[263], stage056[296], stage055[303]}
   );
   gpc1_1 gpc1_1_8786(
      {stage058[238]},
      {stage058[240]}
   );
   gpc3_2 gpc3_2_8787(
      {stage059[321], stage059[322], stage059[323]},
      {stage060[252], stage059[325]}
   );
   gpc2135_5 gpc2135_5_8788(
      {stage060[247], stage060[248], stage060[249], stage060[250], stage060[251]},
      {stage061[281], stage061[282], 1'h0},
      {stage062[259]},
      {stage063[219], stage063[220]},
      {stage064[271], stage063[225], stage062[261], stage061[283], stage060[253]}
   );
   gpc1343_5 gpc1343_5_8789(
      {stage062[260], 1'h0, 1'h0},
      {stage063[221], stage063[222], stage063[223], stage063[224]},
      {stage064[269], stage064[270], 1'h0},
      {stage065[264]},
      {stage066[291], stage065[268], stage064[272], stage063[226], stage062[262]}
   );
   gpc215_4 gpc215_4_8790(
      {stage065[265], stage065[266], stage065[267], 1'h0, 1'h0},
      {stage066[290]},
      {stage067[268], stage067[269]},
      {stage068[287], stage067[270], stage066[292], stage065[269]}
   );
   gpc7_3 gpc7_3_8791(
      {stage068[281], stage068[282], stage068[283], stage068[284], stage068[285], stage068[286], 1'h0},
      {stage070[268], stage069[276], stage068[288]}
   );
   gpc2135_5 gpc2135_5_8792(
      {stage069[272], stage069[273], stage069[274], stage069[275], 1'h0},
      {stage070[265], stage070[266], stage070[267]},
      {stage071[266]},
      {stage072[315], 1'h0},
      {stage073[251], stage072[316], stage071[270], stage070[269], stage069[277]}
   );
   gpc606_5 gpc606_5_8793(
      {stage071[267], stage071[268], stage071[269], 1'h0, 1'h0, 1'h0},
      {stage073[247], stage073[248], stage073[249], stage073[250], 1'h0, 1'h0},
      {stage075[214], stage074[266], stage073[252], stage072[317], stage071[271]}
   );
   gpc135_4 gpc135_4_8794(
      {stage074[262], stage074[263], stage074[264], stage074[265], 1'h0},
      {stage075[212], stage075[213], 1'h0},
      {stage076[218]},
      {stage077[269], stage076[220], stage075[215], stage074[267]}
   );
   gpc1_1 gpc1_1_8795(
      {stage076[219]},
      {stage076[221]}
   );
   gpc7_3 gpc7_3_8796(
      {stage077[263], stage077[264], stage077[265], stage077[266], stage077[267], stage077[268], 1'h0},
      {stage079[263], stage078[238], stage077[270]}
   );
   gpc135_4 gpc135_4_8797(
      {stage078[235], stage078[236], stage078[237], 1'h0, 1'h0},
      {stage079[260], stage079[261], stage079[262]},
      {stage080[266]},
      {stage081[298], stage080[268], stage079[264], stage078[239]}
   );
   gpc1_1 gpc1_1_8798(
      {stage080[267]},
      {stage080[269]}
   );
   gpc615_5 gpc615_5_8799(
      {stage081[293], stage081[294], stage081[295], stage081[296], stage081[297]},
      {stage082[269]},
      {stage083[277], stage083[278], stage083[279], stage083[280], stage083[281], 1'h0},
      {stage085[279], stage084[248], stage083[282], stage082[271], stage081[299]}
   );
   gpc1_1 gpc1_1_8800(
      {stage082[270]},
      {stage082[272]}
   );
   gpc1325_5 gpc1325_5_8801(
      {stage084[243], stage084[244], stage084[245], stage084[246], stage084[247]},
      {stage085[277], stage085[278]},
      {stage086[292], stage086[293], stage086[294]},
      {stage087[242]},
      {stage088[286], stage087[244], stage086[296], stage085[280], stage084[249]}
   );
   gpc1_1 gpc1_1_8802(
      {stage086[295]},
      {stage086[297]}
   );
   gpc1_1 gpc1_1_8803(
      {stage087[243]},
      {stage087[245]}
   );
   gpc606_5 gpc606_5_8804(
      {stage088[282], stage088[283], stage088[284], stage088[285], 1'h0, 1'h0},
      {stage090[253], stage090[254], stage090[255], stage090[256], stage090[257], stage090[258]},
      {stage092[258], stage091[344], stage090[259], stage089[276], stage088[287]}
   );
   gpc3_2 gpc3_2_8805(
      {stage089[273], stage089[274], stage089[275]},
      {stage090[260], stage089[277]}
   );
   gpc135_4 gpc135_4_8806(
      {stage091[339], stage091[340], stage091[341], stage091[342], stage091[343]},
      {stage092[255], stage092[256], stage092[257]},
      {stage093[239]},
      {stage094[250], stage093[241], stage092[259], stage091[345]}
   );
   gpc1_1 gpc1_1_8807(
      {stage093[240]},
      {stage093[242]}
   );
   gpc207_4 gpc207_4_8808(
      {stage094[244], stage094[245], stage094[246], stage094[247], stage094[248], stage094[249], 1'h0},
      {stage096[244], stage096[245]},
      {stage097[233], stage096[247], stage095[230], stage094[251]}
   );
   gpc615_5 gpc615_5_8809(
      {stage095[225], stage095[226], stage095[227], stage095[228], stage095[229]},
      {stage096[246]},
      {stage097[229], stage097[230], stage097[231], stage097[232], 1'h0, 1'h0},
      {stage099[303], stage098[245], stage097[234], stage096[248], stage095[231]}
   );
   gpc1_1 gpc1_1_8810(
      {stage098[244]},
      {stage098[246]}
   );
   gpc7_3 gpc7_3_8811(
      {stage099[296], stage099[297], stage099[298], stage099[299], stage099[300], stage099[301], stage099[302]},
      {stage101[271], stage100[230], stage099[304]}
   );
   gpc1_1 gpc1_1_8812(
      {stage100[229]},
      {stage100[231]}
   );
   gpc1406_5 gpc1406_5_8813(
      {stage101[265], stage101[266], stage101[267], stage101[268], stage101[269], stage101[270]},
      {stage103[255], stage103[256], stage103[257], stage103[258]},
      {stage104[265]},
      {stage105[230], stage104[266], stage103[261], stage102[251], stage101[272]}
   );
   gpc23_3 gpc23_3_8814(
      {stage102[249], stage102[250], 1'h0},
      {stage103[259], stage103[260]},
      {stage104[267], stage103[262], stage102[252]}
   );
   gpc615_5 gpc615_5_8815(
      {stage105[226], stage105[227], stage105[228], stage105[229], 1'h0},
      {stage106[256]},
      {stage107[261], stage107[262], stage107[263], stage107[264], stage107[265], stage107[266]},
      {stage109[236], stage108[264], stage107[267], stage106[260], stage105[231]}
   );
   gpc1406_5 gpc1406_5_8816(
      {stage106[257], stage106[258], stage106[259], 1'h0, 1'h0, 1'h0},
      {stage108[263], 1'h0, 1'h0, 1'h0},
      {stage109[235]},
      {stage110[272], stage109[237], stage108[265], stage107[268], stage106[261]}
   );
   gpc615_5 gpc615_5_8817(
      {stage110[268], stage110[269], stage110[270], stage110[271], 1'h0},
      {stage111[263]},
      {stage112[239], stage112[240], stage112[241], stage112[242], stage112[243], 1'h0},
      {stage114[253], stage113[242], stage112[244], stage111[265], stage110[273]}
   );
   gpc1_1 gpc1_1_8818(
      {stage111[264]},
      {stage111[266]}
   );
   gpc1_1 gpc1_1_8819(
      {stage113[241]},
      {stage113[243]}
   );
   gpc207_4 gpc207_4_8820(
      {stage114[247], stage114[248], stage114[249], stage114[250], stage114[251], stage114[252], 1'h0},
      {stage116[241], stage116[242]},
      {stage117[264], stage116[243], stage115[263], stage114[254]}
   );
   gpc606_5 gpc606_5_8821(
      {stage115[261], stage115[262], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage117[258], stage117[259], stage117[260], stage117[261], stage117[262], stage117[263]},
      {stage119[241], stage118[264], stage117[265], stage116[244], stage115[264]}
   );
   gpc1_1 gpc1_1_8822(
      {stage118[263]},
      {stage118[265]}
   );
   gpc606_5 gpc606_5_8823(
      {stage119[236], stage119[237], stage119[238], stage119[239], stage119[240], 1'h0},
      {stage121[235], stage121[236], stage121[237], stage121[238], stage121[239], stage121[240]},
      {stage123[328], stage122[249], stage121[241], stage120[256], stage119[242]}
   );
   gpc1_1 gpc1_1_8824(
      {stage120[255]},
      {stage120[257]}
   );
   gpc223_4 gpc223_4_8825(
      {stage122[246], stage122[247], stage122[248]},
      {stage123[326], stage123[327]},
      {stage124[236], stage124[237]},
      {stage125[286], stage124[239], stage123[329], stage122[250]}
   );
   gpc1_1 gpc1_1_8826(
      {stage124[238]},
      {stage124[240]}
   );
   gpc23_3 gpc23_3_8827(
      {stage125[283], stage125[284], stage125[285]},
      {stage126[284], stage126[285]},
      {stage127[291], stage126[287], stage125[287]}
   );
   gpc1_1 gpc1_1_8828(
      {stage126[286]},
      {stage126[288]}
   );
   gpc23_3 gpc23_3_8829(
      {stage127[288], stage127[289], stage127[290]},
      {stage128[87], stage128[88]},
      {stage129[86], stage128[90], stage127[292]}
   );
   gpc1_1 gpc1_1_8830(
      {stage128[89]},
      {stage128[91]}
   );
   gpc207_4 gpc207_4_8831(
      {stage129[80], stage129[81], stage129[82], stage129[83], stage129[84], stage129[85], 1'h0},
      {stage131[11], stage131[12]},
      {stage132[7], stage131[16], stage130[20], stage129[87]}
   );
   gpc2135_5 gpc2135_5_8832(
      {stage130[17], stage130[18], stage130[19], 1'h0, 1'h0},
      {stage131[13], stage131[14], stage131[15]},
      {stage132[6]},
      {stage133[3], stage133[4]},
      {stage134[0], stage133[6], stage132[8], stage131[17], stage130[21]}
   );
   gpc1_1 gpc1_1_8833(
      {stage133[5]},
      {stage133[7]}
   );
endmodule

module behavioral_tester();
   reg [127:0] src000;
   reg [127:0] src001;
   reg [127:0] src002;
   reg [127:0] src003;
   reg [127:0] src004;
   reg [127:0] src005;
   reg [127:0] src006;
   reg [127:0] src007;
   reg [127:0] src008;
   reg [127:0] src009;
   reg [127:0] src010;
   reg [127:0] src011;
   reg [127:0] src012;
   reg [127:0] src013;
   reg [127:0] src014;
   reg [127:0] src015;
   reg [127:0] src016;
   reg [127:0] src017;
   reg [127:0] src018;
   reg [127:0] src019;
   reg [127:0] src020;
   reg [127:0] src021;
   reg [127:0] src022;
   reg [127:0] src023;
   reg [127:0] src024;
   reg [127:0] src025;
   reg [127:0] src026;
   reg [127:0] src027;
   reg [127:0] src028;
   reg [127:0] src029;
   reg [127:0] src030;
   reg [127:0] src031;
   reg [127:0] src032;
   reg [127:0] src033;
   reg [127:0] src034;
   reg [127:0] src035;
   reg [127:0] src036;
   reg [127:0] src037;
   reg [127:0] src038;
   reg [127:0] src039;
   reg [127:0] src040;
   reg [127:0] src041;
   reg [127:0] src042;
   reg [127:0] src043;
   reg [127:0] src044;
   reg [127:0] src045;
   reg [127:0] src046;
   reg [127:0] src047;
   reg [127:0] src048;
   reg [127:0] src049;
   reg [127:0] src050;
   reg [127:0] src051;
   reg [127:0] src052;
   reg [127:0] src053;
   reg [127:0] src054;
   reg [127:0] src055;
   reg [127:0] src056;
   reg [127:0] src057;
   reg [127:0] src058;
   reg [127:0] src059;
   reg [127:0] src060;
   reg [127:0] src061;
   reg [127:0] src062;
   reg [127:0] src063;
   reg [127:0] src064;
   reg [127:0] src065;
   reg [127:0] src066;
   reg [127:0] src067;
   reg [127:0] src068;
   reg [127:0] src069;
   reg [127:0] src070;
   reg [127:0] src071;
   reg [127:0] src072;
   reg [127:0] src073;
   reg [127:0] src074;
   reg [127:0] src075;
   reg [127:0] src076;
   reg [127:0] src077;
   reg [127:0] src078;
   reg [127:0] src079;
   reg [127:0] src080;
   reg [127:0] src081;
   reg [127:0] src082;
   reg [127:0] src083;
   reg [127:0] src084;
   reg [127:0] src085;
   reg [127:0] src086;
   reg [127:0] src087;
   reg [127:0] src088;
   reg [127:0] src089;
   reg [127:0] src090;
   reg [127:0] src091;
   reg [127:0] src092;
   reg [127:0] src093;
   reg [127:0] src094;
   reg [127:0] src095;
   reg [127:0] src096;
   reg [127:0] src097;
   reg [127:0] src098;
   reg [127:0] src099;
   reg [127:0] src100;
   reg [127:0] src101;
   reg [127:0] src102;
   reg [127:0] src103;
   reg [127:0] src104;
   reg [127:0] src105;
   reg [127:0] src106;
   reg [127:0] src107;
   reg [127:0] src108;
   reg [127:0] src109;
   reg [127:0] src110;
   reg [127:0] src111;
   reg [127:0] src112;
   reg [127:0] src113;
   reg [127:0] src114;
   reg [127:0] src115;
   reg [127:0] src116;
   reg [127:0] src117;
   reg [127:0] src118;
   reg [127:0] src119;
   reg [127:0] src120;
   reg [127:0] src121;
   reg [127:0] src122;
   reg [127:0] src123;
   reg [127:0] src124;
   reg [127:0] src125;
   reg [127:0] src126;
   reg [127:0] src127;
   wire [1:0] dst000;
   wire [1:0] dst001;
   wire [1:0] dst002;
   wire [0:0] dst003;
   wire [0:0] dst004;
   wire [1:0] dst005;
   wire [0:0] dst006;
   wire [1:0] dst007;
   wire [1:0] dst008;
   wire [1:0] dst009;
   wire [1:0] dst010;
   wire [1:0] dst011;
   wire [1:0] dst012;
   wire [0:0] dst013;
   wire [1:0] dst014;
   wire [1:0] dst015;
   wire [1:0] dst016;
   wire [1:0] dst017;
   wire [1:0] dst018;
   wire [1:0] dst019;
   wire [1:0] dst020;
   wire [1:0] dst021;
   wire [1:0] dst022;
   wire [1:0] dst023;
   wire [1:0] dst024;
   wire [1:0] dst025;
   wire [1:0] dst026;
   wire [1:0] dst027;
   wire [1:0] dst028;
   wire [1:0] dst029;
   wire [1:0] dst030;
   wire [1:0] dst031;
   wire [1:0] dst032;
   wire [1:0] dst033;
   wire [1:0] dst034;
   wire [1:0] dst035;
   wire [1:0] dst036;
   wire [1:0] dst037;
   wire [0:0] dst038;
   wire [0:0] dst039;
   wire [1:0] dst040;
   wire [1:0] dst041;
   wire [1:0] dst042;
   wire [1:0] dst043;
   wire [1:0] dst044;
   wire [1:0] dst045;
   wire [1:0] dst046;
   wire [1:0] dst047;
   wire [1:0] dst048;
   wire [1:0] dst049;
   wire [1:0] dst050;
   wire [1:0] dst051;
   wire [1:0] dst052;
   wire [1:0] dst053;
   wire [1:0] dst054;
   wire [1:0] dst055;
   wire [1:0] dst056;
   wire [1:0] dst057;
   wire [1:0] dst058;
   wire [1:0] dst059;
   wire [1:0] dst060;
   wire [0:0] dst061;
   wire [1:0] dst062;
   wire [1:0] dst063;
   wire [1:0] dst064;
   wire [1:0] dst065;
   wire [1:0] dst066;
   wire [0:0] dst067;
   wire [1:0] dst068;
   wire [1:0] dst069;
   wire [1:0] dst070;
   wire [1:0] dst071;
   wire [1:0] dst072;
   wire [1:0] dst073;
   wire [1:0] dst074;
   wire [1:0] dst075;
   wire [1:0] dst076;
   wire [1:0] dst077;
   wire [1:0] dst078;
   wire [1:0] dst079;
   wire [1:0] dst080;
   wire [1:0] dst081;
   wire [1:0] dst082;
   wire [0:0] dst083;
   wire [1:0] dst084;
   wire [1:0] dst085;
   wire [1:0] dst086;
   wire [1:0] dst087;
   wire [1:0] dst088;
   wire [1:0] dst089;
   wire [1:0] dst090;
   wire [1:0] dst091;
   wire [1:0] dst092;
   wire [1:0] dst093;
   wire [1:0] dst094;
   wire [1:0] dst095;
   wire [1:0] dst096;
   wire [1:0] dst097;
   wire [1:0] dst098;
   wire [1:0] dst099;
   wire [1:0] dst100;
   wire [1:0] dst101;
   wire [1:0] dst102;
   wire [1:0] dst103;
   wire [1:0] dst104;
   wire [1:0] dst105;
   wire [1:0] dst106;
   wire [1:0] dst107;
   wire [1:0] dst108;
   wire [1:0] dst109;
   wire [1:0] dst110;
   wire [1:0] dst111;
   wire [0:0] dst112;
   wire [1:0] dst113;
   wire [1:0] dst114;
   wire [1:0] dst115;
   wire [1:0] dst116;
   wire [1:0] dst117;
   wire [1:0] dst118;
   wire [1:0] dst119;
   wire [1:0] dst120;
   wire [0:0] dst121;
   wire [1:0] dst122;
   wire [1:0] dst123;
   wire [1:0] dst124;
   wire [1:0] dst125;
   wire [1:0] dst126;
   wire [1:0] dst127;
   wire [1:0] dst128;
   wire [1:0] dst129;
   wire [1:0] dst130;
   wire [1:0] dst131;
   wire [1:0] dst132;
   wire [1:0] dst133;
   wire [0:0] dst134;
   wire [135:0] srcsum;
   wire [135:0] dstsum;
   wire test;
   assign srcsum =
      (src000[0] << 0) +
      (src000[1] << 0) +
      (src000[2] << 0) +
      (src000[3] << 0) +
      (src000[4] << 0) +
      (src000[5] << 0) +
      (src000[6] << 0) +
      (src000[7] << 0) +
      (src000[8] << 0) +
      (src000[9] << 0) +
      (src000[10] << 0) +
      (src000[11] << 0) +
      (src000[12] << 0) +
      (src000[13] << 0) +
      (src000[14] << 0) +
      (src000[15] << 0) +
      (src000[16] << 0) +
      (src000[17] << 0) +
      (src000[18] << 0) +
      (src000[19] << 0) +
      (src000[20] << 0) +
      (src000[21] << 0) +
      (src000[22] << 0) +
      (src000[23] << 0) +
      (src000[24] << 0) +
      (src000[25] << 0) +
      (src000[26] << 0) +
      (src000[27] << 0) +
      (src000[28] << 0) +
      (src000[29] << 0) +
      (src000[30] << 0) +
      (src000[31] << 0) +
      (src000[32] << 0) +
      (src000[33] << 0) +
      (src000[34] << 0) +
      (src000[35] << 0) +
      (src000[36] << 0) +
      (src000[37] << 0) +
      (src000[38] << 0) +
      (src000[39] << 0) +
      (src000[40] << 0) +
      (src000[41] << 0) +
      (src000[42] << 0) +
      (src000[43] << 0) +
      (src000[44] << 0) +
      (src000[45] << 0) +
      (src000[46] << 0) +
      (src000[47] << 0) +
      (src000[48] << 0) +
      (src000[49] << 0) +
      (src000[50] << 0) +
      (src000[51] << 0) +
      (src000[52] << 0) +
      (src000[53] << 0) +
      (src000[54] << 0) +
      (src000[55] << 0) +
      (src000[56] << 0) +
      (src000[57] << 0) +
      (src000[58] << 0) +
      (src000[59] << 0) +
      (src000[60] << 0) +
      (src000[61] << 0) +
      (src000[62] << 0) +
      (src000[63] << 0) +
      (src000[64] << 0) +
      (src000[65] << 0) +
      (src000[66] << 0) +
      (src000[67] << 0) +
      (src000[68] << 0) +
      (src000[69] << 0) +
      (src000[70] << 0) +
      (src000[71] << 0) +
      (src000[72] << 0) +
      (src000[73] << 0) +
      (src000[74] << 0) +
      (src000[75] << 0) +
      (src000[76] << 0) +
      (src000[77] << 0) +
      (src000[78] << 0) +
      (src000[79] << 0) +
      (src000[80] << 0) +
      (src000[81] << 0) +
      (src000[82] << 0) +
      (src000[83] << 0) +
      (src000[84] << 0) +
      (src000[85] << 0) +
      (src000[86] << 0) +
      (src000[87] << 0) +
      (src000[88] << 0) +
      (src000[89] << 0) +
      (src000[90] << 0) +
      (src000[91] << 0) +
      (src000[92] << 0) +
      (src000[93] << 0) +
      (src000[94] << 0) +
      (src000[95] << 0) +
      (src000[96] << 0) +
      (src000[97] << 0) +
      (src000[98] << 0) +
      (src000[99] << 0) +
      (src000[100] << 0) +
      (src000[101] << 0) +
      (src000[102] << 0) +
      (src000[103] << 0) +
      (src000[104] << 0) +
      (src000[105] << 0) +
      (src000[106] << 0) +
      (src000[107] << 0) +
      (src000[108] << 0) +
      (src000[109] << 0) +
      (src000[110] << 0) +
      (src000[111] << 0) +
      (src000[112] << 0) +
      (src000[113] << 0) +
      (src000[114] << 0) +
      (src000[115] << 0) +
      (src000[116] << 0) +
      (src000[117] << 0) +
      (src000[118] << 0) +
      (src000[119] << 0) +
      (src000[120] << 0) +
      (src000[121] << 0) +
      (src000[122] << 0) +
      (src000[123] << 0) +
      (src000[124] << 0) +
      (src000[125] << 0) +
      (src000[126] << 0) +
      (src000[127] << 0) +
      (src001[0] << 1) +
      (src001[1] << 1) +
      (src001[2] << 1) +
      (src001[3] << 1) +
      (src001[4] << 1) +
      (src001[5] << 1) +
      (src001[6] << 1) +
      (src001[7] << 1) +
      (src001[8] << 1) +
      (src001[9] << 1) +
      (src001[10] << 1) +
      (src001[11] << 1) +
      (src001[12] << 1) +
      (src001[13] << 1) +
      (src001[14] << 1) +
      (src001[15] << 1) +
      (src001[16] << 1) +
      (src001[17] << 1) +
      (src001[18] << 1) +
      (src001[19] << 1) +
      (src001[20] << 1) +
      (src001[21] << 1) +
      (src001[22] << 1) +
      (src001[23] << 1) +
      (src001[24] << 1) +
      (src001[25] << 1) +
      (src001[26] << 1) +
      (src001[27] << 1) +
      (src001[28] << 1) +
      (src001[29] << 1) +
      (src001[30] << 1) +
      (src001[31] << 1) +
      (src001[32] << 1) +
      (src001[33] << 1) +
      (src001[34] << 1) +
      (src001[35] << 1) +
      (src001[36] << 1) +
      (src001[37] << 1) +
      (src001[38] << 1) +
      (src001[39] << 1) +
      (src001[40] << 1) +
      (src001[41] << 1) +
      (src001[42] << 1) +
      (src001[43] << 1) +
      (src001[44] << 1) +
      (src001[45] << 1) +
      (src001[46] << 1) +
      (src001[47] << 1) +
      (src001[48] << 1) +
      (src001[49] << 1) +
      (src001[50] << 1) +
      (src001[51] << 1) +
      (src001[52] << 1) +
      (src001[53] << 1) +
      (src001[54] << 1) +
      (src001[55] << 1) +
      (src001[56] << 1) +
      (src001[57] << 1) +
      (src001[58] << 1) +
      (src001[59] << 1) +
      (src001[60] << 1) +
      (src001[61] << 1) +
      (src001[62] << 1) +
      (src001[63] << 1) +
      (src001[64] << 1) +
      (src001[65] << 1) +
      (src001[66] << 1) +
      (src001[67] << 1) +
      (src001[68] << 1) +
      (src001[69] << 1) +
      (src001[70] << 1) +
      (src001[71] << 1) +
      (src001[72] << 1) +
      (src001[73] << 1) +
      (src001[74] << 1) +
      (src001[75] << 1) +
      (src001[76] << 1) +
      (src001[77] << 1) +
      (src001[78] << 1) +
      (src001[79] << 1) +
      (src001[80] << 1) +
      (src001[81] << 1) +
      (src001[82] << 1) +
      (src001[83] << 1) +
      (src001[84] << 1) +
      (src001[85] << 1) +
      (src001[86] << 1) +
      (src001[87] << 1) +
      (src001[88] << 1) +
      (src001[89] << 1) +
      (src001[90] << 1) +
      (src001[91] << 1) +
      (src001[92] << 1) +
      (src001[93] << 1) +
      (src001[94] << 1) +
      (src001[95] << 1) +
      (src001[96] << 1) +
      (src001[97] << 1) +
      (src001[98] << 1) +
      (src001[99] << 1) +
      (src001[100] << 1) +
      (src001[101] << 1) +
      (src001[102] << 1) +
      (src001[103] << 1) +
      (src001[104] << 1) +
      (src001[105] << 1) +
      (src001[106] << 1) +
      (src001[107] << 1) +
      (src001[108] << 1) +
      (src001[109] << 1) +
      (src001[110] << 1) +
      (src001[111] << 1) +
      (src001[112] << 1) +
      (src001[113] << 1) +
      (src001[114] << 1) +
      (src001[115] << 1) +
      (src001[116] << 1) +
      (src001[117] << 1) +
      (src001[118] << 1) +
      (src001[119] << 1) +
      (src001[120] << 1) +
      (src001[121] << 1) +
      (src001[122] << 1) +
      (src001[123] << 1) +
      (src001[124] << 1) +
      (src001[125] << 1) +
      (src001[126] << 1) +
      (src001[127] << 1) +
      (src002[0] << 2) +
      (src002[1] << 2) +
      (src002[2] << 2) +
      (src002[3] << 2) +
      (src002[4] << 2) +
      (src002[5] << 2) +
      (src002[6] << 2) +
      (src002[7] << 2) +
      (src002[8] << 2) +
      (src002[9] << 2) +
      (src002[10] << 2) +
      (src002[11] << 2) +
      (src002[12] << 2) +
      (src002[13] << 2) +
      (src002[14] << 2) +
      (src002[15] << 2) +
      (src002[16] << 2) +
      (src002[17] << 2) +
      (src002[18] << 2) +
      (src002[19] << 2) +
      (src002[20] << 2) +
      (src002[21] << 2) +
      (src002[22] << 2) +
      (src002[23] << 2) +
      (src002[24] << 2) +
      (src002[25] << 2) +
      (src002[26] << 2) +
      (src002[27] << 2) +
      (src002[28] << 2) +
      (src002[29] << 2) +
      (src002[30] << 2) +
      (src002[31] << 2) +
      (src002[32] << 2) +
      (src002[33] << 2) +
      (src002[34] << 2) +
      (src002[35] << 2) +
      (src002[36] << 2) +
      (src002[37] << 2) +
      (src002[38] << 2) +
      (src002[39] << 2) +
      (src002[40] << 2) +
      (src002[41] << 2) +
      (src002[42] << 2) +
      (src002[43] << 2) +
      (src002[44] << 2) +
      (src002[45] << 2) +
      (src002[46] << 2) +
      (src002[47] << 2) +
      (src002[48] << 2) +
      (src002[49] << 2) +
      (src002[50] << 2) +
      (src002[51] << 2) +
      (src002[52] << 2) +
      (src002[53] << 2) +
      (src002[54] << 2) +
      (src002[55] << 2) +
      (src002[56] << 2) +
      (src002[57] << 2) +
      (src002[58] << 2) +
      (src002[59] << 2) +
      (src002[60] << 2) +
      (src002[61] << 2) +
      (src002[62] << 2) +
      (src002[63] << 2) +
      (src002[64] << 2) +
      (src002[65] << 2) +
      (src002[66] << 2) +
      (src002[67] << 2) +
      (src002[68] << 2) +
      (src002[69] << 2) +
      (src002[70] << 2) +
      (src002[71] << 2) +
      (src002[72] << 2) +
      (src002[73] << 2) +
      (src002[74] << 2) +
      (src002[75] << 2) +
      (src002[76] << 2) +
      (src002[77] << 2) +
      (src002[78] << 2) +
      (src002[79] << 2) +
      (src002[80] << 2) +
      (src002[81] << 2) +
      (src002[82] << 2) +
      (src002[83] << 2) +
      (src002[84] << 2) +
      (src002[85] << 2) +
      (src002[86] << 2) +
      (src002[87] << 2) +
      (src002[88] << 2) +
      (src002[89] << 2) +
      (src002[90] << 2) +
      (src002[91] << 2) +
      (src002[92] << 2) +
      (src002[93] << 2) +
      (src002[94] << 2) +
      (src002[95] << 2) +
      (src002[96] << 2) +
      (src002[97] << 2) +
      (src002[98] << 2) +
      (src002[99] << 2) +
      (src002[100] << 2) +
      (src002[101] << 2) +
      (src002[102] << 2) +
      (src002[103] << 2) +
      (src002[104] << 2) +
      (src002[105] << 2) +
      (src002[106] << 2) +
      (src002[107] << 2) +
      (src002[108] << 2) +
      (src002[109] << 2) +
      (src002[110] << 2) +
      (src002[111] << 2) +
      (src002[112] << 2) +
      (src002[113] << 2) +
      (src002[114] << 2) +
      (src002[115] << 2) +
      (src002[116] << 2) +
      (src002[117] << 2) +
      (src002[118] << 2) +
      (src002[119] << 2) +
      (src002[120] << 2) +
      (src002[121] << 2) +
      (src002[122] << 2) +
      (src002[123] << 2) +
      (src002[124] << 2) +
      (src002[125] << 2) +
      (src002[126] << 2) +
      (src002[127] << 2) +
      (src003[0] << 3) +
      (src003[1] << 3) +
      (src003[2] << 3) +
      (src003[3] << 3) +
      (src003[4] << 3) +
      (src003[5] << 3) +
      (src003[6] << 3) +
      (src003[7] << 3) +
      (src003[8] << 3) +
      (src003[9] << 3) +
      (src003[10] << 3) +
      (src003[11] << 3) +
      (src003[12] << 3) +
      (src003[13] << 3) +
      (src003[14] << 3) +
      (src003[15] << 3) +
      (src003[16] << 3) +
      (src003[17] << 3) +
      (src003[18] << 3) +
      (src003[19] << 3) +
      (src003[20] << 3) +
      (src003[21] << 3) +
      (src003[22] << 3) +
      (src003[23] << 3) +
      (src003[24] << 3) +
      (src003[25] << 3) +
      (src003[26] << 3) +
      (src003[27] << 3) +
      (src003[28] << 3) +
      (src003[29] << 3) +
      (src003[30] << 3) +
      (src003[31] << 3) +
      (src003[32] << 3) +
      (src003[33] << 3) +
      (src003[34] << 3) +
      (src003[35] << 3) +
      (src003[36] << 3) +
      (src003[37] << 3) +
      (src003[38] << 3) +
      (src003[39] << 3) +
      (src003[40] << 3) +
      (src003[41] << 3) +
      (src003[42] << 3) +
      (src003[43] << 3) +
      (src003[44] << 3) +
      (src003[45] << 3) +
      (src003[46] << 3) +
      (src003[47] << 3) +
      (src003[48] << 3) +
      (src003[49] << 3) +
      (src003[50] << 3) +
      (src003[51] << 3) +
      (src003[52] << 3) +
      (src003[53] << 3) +
      (src003[54] << 3) +
      (src003[55] << 3) +
      (src003[56] << 3) +
      (src003[57] << 3) +
      (src003[58] << 3) +
      (src003[59] << 3) +
      (src003[60] << 3) +
      (src003[61] << 3) +
      (src003[62] << 3) +
      (src003[63] << 3) +
      (src003[64] << 3) +
      (src003[65] << 3) +
      (src003[66] << 3) +
      (src003[67] << 3) +
      (src003[68] << 3) +
      (src003[69] << 3) +
      (src003[70] << 3) +
      (src003[71] << 3) +
      (src003[72] << 3) +
      (src003[73] << 3) +
      (src003[74] << 3) +
      (src003[75] << 3) +
      (src003[76] << 3) +
      (src003[77] << 3) +
      (src003[78] << 3) +
      (src003[79] << 3) +
      (src003[80] << 3) +
      (src003[81] << 3) +
      (src003[82] << 3) +
      (src003[83] << 3) +
      (src003[84] << 3) +
      (src003[85] << 3) +
      (src003[86] << 3) +
      (src003[87] << 3) +
      (src003[88] << 3) +
      (src003[89] << 3) +
      (src003[90] << 3) +
      (src003[91] << 3) +
      (src003[92] << 3) +
      (src003[93] << 3) +
      (src003[94] << 3) +
      (src003[95] << 3) +
      (src003[96] << 3) +
      (src003[97] << 3) +
      (src003[98] << 3) +
      (src003[99] << 3) +
      (src003[100] << 3) +
      (src003[101] << 3) +
      (src003[102] << 3) +
      (src003[103] << 3) +
      (src003[104] << 3) +
      (src003[105] << 3) +
      (src003[106] << 3) +
      (src003[107] << 3) +
      (src003[108] << 3) +
      (src003[109] << 3) +
      (src003[110] << 3) +
      (src003[111] << 3) +
      (src003[112] << 3) +
      (src003[113] << 3) +
      (src003[114] << 3) +
      (src003[115] << 3) +
      (src003[116] << 3) +
      (src003[117] << 3) +
      (src003[118] << 3) +
      (src003[119] << 3) +
      (src003[120] << 3) +
      (src003[121] << 3) +
      (src003[122] << 3) +
      (src003[123] << 3) +
      (src003[124] << 3) +
      (src003[125] << 3) +
      (src003[126] << 3) +
      (src003[127] << 3) +
      (src004[0] << 4) +
      (src004[1] << 4) +
      (src004[2] << 4) +
      (src004[3] << 4) +
      (src004[4] << 4) +
      (src004[5] << 4) +
      (src004[6] << 4) +
      (src004[7] << 4) +
      (src004[8] << 4) +
      (src004[9] << 4) +
      (src004[10] << 4) +
      (src004[11] << 4) +
      (src004[12] << 4) +
      (src004[13] << 4) +
      (src004[14] << 4) +
      (src004[15] << 4) +
      (src004[16] << 4) +
      (src004[17] << 4) +
      (src004[18] << 4) +
      (src004[19] << 4) +
      (src004[20] << 4) +
      (src004[21] << 4) +
      (src004[22] << 4) +
      (src004[23] << 4) +
      (src004[24] << 4) +
      (src004[25] << 4) +
      (src004[26] << 4) +
      (src004[27] << 4) +
      (src004[28] << 4) +
      (src004[29] << 4) +
      (src004[30] << 4) +
      (src004[31] << 4) +
      (src004[32] << 4) +
      (src004[33] << 4) +
      (src004[34] << 4) +
      (src004[35] << 4) +
      (src004[36] << 4) +
      (src004[37] << 4) +
      (src004[38] << 4) +
      (src004[39] << 4) +
      (src004[40] << 4) +
      (src004[41] << 4) +
      (src004[42] << 4) +
      (src004[43] << 4) +
      (src004[44] << 4) +
      (src004[45] << 4) +
      (src004[46] << 4) +
      (src004[47] << 4) +
      (src004[48] << 4) +
      (src004[49] << 4) +
      (src004[50] << 4) +
      (src004[51] << 4) +
      (src004[52] << 4) +
      (src004[53] << 4) +
      (src004[54] << 4) +
      (src004[55] << 4) +
      (src004[56] << 4) +
      (src004[57] << 4) +
      (src004[58] << 4) +
      (src004[59] << 4) +
      (src004[60] << 4) +
      (src004[61] << 4) +
      (src004[62] << 4) +
      (src004[63] << 4) +
      (src004[64] << 4) +
      (src004[65] << 4) +
      (src004[66] << 4) +
      (src004[67] << 4) +
      (src004[68] << 4) +
      (src004[69] << 4) +
      (src004[70] << 4) +
      (src004[71] << 4) +
      (src004[72] << 4) +
      (src004[73] << 4) +
      (src004[74] << 4) +
      (src004[75] << 4) +
      (src004[76] << 4) +
      (src004[77] << 4) +
      (src004[78] << 4) +
      (src004[79] << 4) +
      (src004[80] << 4) +
      (src004[81] << 4) +
      (src004[82] << 4) +
      (src004[83] << 4) +
      (src004[84] << 4) +
      (src004[85] << 4) +
      (src004[86] << 4) +
      (src004[87] << 4) +
      (src004[88] << 4) +
      (src004[89] << 4) +
      (src004[90] << 4) +
      (src004[91] << 4) +
      (src004[92] << 4) +
      (src004[93] << 4) +
      (src004[94] << 4) +
      (src004[95] << 4) +
      (src004[96] << 4) +
      (src004[97] << 4) +
      (src004[98] << 4) +
      (src004[99] << 4) +
      (src004[100] << 4) +
      (src004[101] << 4) +
      (src004[102] << 4) +
      (src004[103] << 4) +
      (src004[104] << 4) +
      (src004[105] << 4) +
      (src004[106] << 4) +
      (src004[107] << 4) +
      (src004[108] << 4) +
      (src004[109] << 4) +
      (src004[110] << 4) +
      (src004[111] << 4) +
      (src004[112] << 4) +
      (src004[113] << 4) +
      (src004[114] << 4) +
      (src004[115] << 4) +
      (src004[116] << 4) +
      (src004[117] << 4) +
      (src004[118] << 4) +
      (src004[119] << 4) +
      (src004[120] << 4) +
      (src004[121] << 4) +
      (src004[122] << 4) +
      (src004[123] << 4) +
      (src004[124] << 4) +
      (src004[125] << 4) +
      (src004[126] << 4) +
      (src004[127] << 4) +
      (src005[0] << 5) +
      (src005[1] << 5) +
      (src005[2] << 5) +
      (src005[3] << 5) +
      (src005[4] << 5) +
      (src005[5] << 5) +
      (src005[6] << 5) +
      (src005[7] << 5) +
      (src005[8] << 5) +
      (src005[9] << 5) +
      (src005[10] << 5) +
      (src005[11] << 5) +
      (src005[12] << 5) +
      (src005[13] << 5) +
      (src005[14] << 5) +
      (src005[15] << 5) +
      (src005[16] << 5) +
      (src005[17] << 5) +
      (src005[18] << 5) +
      (src005[19] << 5) +
      (src005[20] << 5) +
      (src005[21] << 5) +
      (src005[22] << 5) +
      (src005[23] << 5) +
      (src005[24] << 5) +
      (src005[25] << 5) +
      (src005[26] << 5) +
      (src005[27] << 5) +
      (src005[28] << 5) +
      (src005[29] << 5) +
      (src005[30] << 5) +
      (src005[31] << 5) +
      (src005[32] << 5) +
      (src005[33] << 5) +
      (src005[34] << 5) +
      (src005[35] << 5) +
      (src005[36] << 5) +
      (src005[37] << 5) +
      (src005[38] << 5) +
      (src005[39] << 5) +
      (src005[40] << 5) +
      (src005[41] << 5) +
      (src005[42] << 5) +
      (src005[43] << 5) +
      (src005[44] << 5) +
      (src005[45] << 5) +
      (src005[46] << 5) +
      (src005[47] << 5) +
      (src005[48] << 5) +
      (src005[49] << 5) +
      (src005[50] << 5) +
      (src005[51] << 5) +
      (src005[52] << 5) +
      (src005[53] << 5) +
      (src005[54] << 5) +
      (src005[55] << 5) +
      (src005[56] << 5) +
      (src005[57] << 5) +
      (src005[58] << 5) +
      (src005[59] << 5) +
      (src005[60] << 5) +
      (src005[61] << 5) +
      (src005[62] << 5) +
      (src005[63] << 5) +
      (src005[64] << 5) +
      (src005[65] << 5) +
      (src005[66] << 5) +
      (src005[67] << 5) +
      (src005[68] << 5) +
      (src005[69] << 5) +
      (src005[70] << 5) +
      (src005[71] << 5) +
      (src005[72] << 5) +
      (src005[73] << 5) +
      (src005[74] << 5) +
      (src005[75] << 5) +
      (src005[76] << 5) +
      (src005[77] << 5) +
      (src005[78] << 5) +
      (src005[79] << 5) +
      (src005[80] << 5) +
      (src005[81] << 5) +
      (src005[82] << 5) +
      (src005[83] << 5) +
      (src005[84] << 5) +
      (src005[85] << 5) +
      (src005[86] << 5) +
      (src005[87] << 5) +
      (src005[88] << 5) +
      (src005[89] << 5) +
      (src005[90] << 5) +
      (src005[91] << 5) +
      (src005[92] << 5) +
      (src005[93] << 5) +
      (src005[94] << 5) +
      (src005[95] << 5) +
      (src005[96] << 5) +
      (src005[97] << 5) +
      (src005[98] << 5) +
      (src005[99] << 5) +
      (src005[100] << 5) +
      (src005[101] << 5) +
      (src005[102] << 5) +
      (src005[103] << 5) +
      (src005[104] << 5) +
      (src005[105] << 5) +
      (src005[106] << 5) +
      (src005[107] << 5) +
      (src005[108] << 5) +
      (src005[109] << 5) +
      (src005[110] << 5) +
      (src005[111] << 5) +
      (src005[112] << 5) +
      (src005[113] << 5) +
      (src005[114] << 5) +
      (src005[115] << 5) +
      (src005[116] << 5) +
      (src005[117] << 5) +
      (src005[118] << 5) +
      (src005[119] << 5) +
      (src005[120] << 5) +
      (src005[121] << 5) +
      (src005[122] << 5) +
      (src005[123] << 5) +
      (src005[124] << 5) +
      (src005[125] << 5) +
      (src005[126] << 5) +
      (src005[127] << 5) +
      (src006[0] << 6) +
      (src006[1] << 6) +
      (src006[2] << 6) +
      (src006[3] << 6) +
      (src006[4] << 6) +
      (src006[5] << 6) +
      (src006[6] << 6) +
      (src006[7] << 6) +
      (src006[8] << 6) +
      (src006[9] << 6) +
      (src006[10] << 6) +
      (src006[11] << 6) +
      (src006[12] << 6) +
      (src006[13] << 6) +
      (src006[14] << 6) +
      (src006[15] << 6) +
      (src006[16] << 6) +
      (src006[17] << 6) +
      (src006[18] << 6) +
      (src006[19] << 6) +
      (src006[20] << 6) +
      (src006[21] << 6) +
      (src006[22] << 6) +
      (src006[23] << 6) +
      (src006[24] << 6) +
      (src006[25] << 6) +
      (src006[26] << 6) +
      (src006[27] << 6) +
      (src006[28] << 6) +
      (src006[29] << 6) +
      (src006[30] << 6) +
      (src006[31] << 6) +
      (src006[32] << 6) +
      (src006[33] << 6) +
      (src006[34] << 6) +
      (src006[35] << 6) +
      (src006[36] << 6) +
      (src006[37] << 6) +
      (src006[38] << 6) +
      (src006[39] << 6) +
      (src006[40] << 6) +
      (src006[41] << 6) +
      (src006[42] << 6) +
      (src006[43] << 6) +
      (src006[44] << 6) +
      (src006[45] << 6) +
      (src006[46] << 6) +
      (src006[47] << 6) +
      (src006[48] << 6) +
      (src006[49] << 6) +
      (src006[50] << 6) +
      (src006[51] << 6) +
      (src006[52] << 6) +
      (src006[53] << 6) +
      (src006[54] << 6) +
      (src006[55] << 6) +
      (src006[56] << 6) +
      (src006[57] << 6) +
      (src006[58] << 6) +
      (src006[59] << 6) +
      (src006[60] << 6) +
      (src006[61] << 6) +
      (src006[62] << 6) +
      (src006[63] << 6) +
      (src006[64] << 6) +
      (src006[65] << 6) +
      (src006[66] << 6) +
      (src006[67] << 6) +
      (src006[68] << 6) +
      (src006[69] << 6) +
      (src006[70] << 6) +
      (src006[71] << 6) +
      (src006[72] << 6) +
      (src006[73] << 6) +
      (src006[74] << 6) +
      (src006[75] << 6) +
      (src006[76] << 6) +
      (src006[77] << 6) +
      (src006[78] << 6) +
      (src006[79] << 6) +
      (src006[80] << 6) +
      (src006[81] << 6) +
      (src006[82] << 6) +
      (src006[83] << 6) +
      (src006[84] << 6) +
      (src006[85] << 6) +
      (src006[86] << 6) +
      (src006[87] << 6) +
      (src006[88] << 6) +
      (src006[89] << 6) +
      (src006[90] << 6) +
      (src006[91] << 6) +
      (src006[92] << 6) +
      (src006[93] << 6) +
      (src006[94] << 6) +
      (src006[95] << 6) +
      (src006[96] << 6) +
      (src006[97] << 6) +
      (src006[98] << 6) +
      (src006[99] << 6) +
      (src006[100] << 6) +
      (src006[101] << 6) +
      (src006[102] << 6) +
      (src006[103] << 6) +
      (src006[104] << 6) +
      (src006[105] << 6) +
      (src006[106] << 6) +
      (src006[107] << 6) +
      (src006[108] << 6) +
      (src006[109] << 6) +
      (src006[110] << 6) +
      (src006[111] << 6) +
      (src006[112] << 6) +
      (src006[113] << 6) +
      (src006[114] << 6) +
      (src006[115] << 6) +
      (src006[116] << 6) +
      (src006[117] << 6) +
      (src006[118] << 6) +
      (src006[119] << 6) +
      (src006[120] << 6) +
      (src006[121] << 6) +
      (src006[122] << 6) +
      (src006[123] << 6) +
      (src006[124] << 6) +
      (src006[125] << 6) +
      (src006[126] << 6) +
      (src006[127] << 6) +
      (src007[0] << 7) +
      (src007[1] << 7) +
      (src007[2] << 7) +
      (src007[3] << 7) +
      (src007[4] << 7) +
      (src007[5] << 7) +
      (src007[6] << 7) +
      (src007[7] << 7) +
      (src007[8] << 7) +
      (src007[9] << 7) +
      (src007[10] << 7) +
      (src007[11] << 7) +
      (src007[12] << 7) +
      (src007[13] << 7) +
      (src007[14] << 7) +
      (src007[15] << 7) +
      (src007[16] << 7) +
      (src007[17] << 7) +
      (src007[18] << 7) +
      (src007[19] << 7) +
      (src007[20] << 7) +
      (src007[21] << 7) +
      (src007[22] << 7) +
      (src007[23] << 7) +
      (src007[24] << 7) +
      (src007[25] << 7) +
      (src007[26] << 7) +
      (src007[27] << 7) +
      (src007[28] << 7) +
      (src007[29] << 7) +
      (src007[30] << 7) +
      (src007[31] << 7) +
      (src007[32] << 7) +
      (src007[33] << 7) +
      (src007[34] << 7) +
      (src007[35] << 7) +
      (src007[36] << 7) +
      (src007[37] << 7) +
      (src007[38] << 7) +
      (src007[39] << 7) +
      (src007[40] << 7) +
      (src007[41] << 7) +
      (src007[42] << 7) +
      (src007[43] << 7) +
      (src007[44] << 7) +
      (src007[45] << 7) +
      (src007[46] << 7) +
      (src007[47] << 7) +
      (src007[48] << 7) +
      (src007[49] << 7) +
      (src007[50] << 7) +
      (src007[51] << 7) +
      (src007[52] << 7) +
      (src007[53] << 7) +
      (src007[54] << 7) +
      (src007[55] << 7) +
      (src007[56] << 7) +
      (src007[57] << 7) +
      (src007[58] << 7) +
      (src007[59] << 7) +
      (src007[60] << 7) +
      (src007[61] << 7) +
      (src007[62] << 7) +
      (src007[63] << 7) +
      (src007[64] << 7) +
      (src007[65] << 7) +
      (src007[66] << 7) +
      (src007[67] << 7) +
      (src007[68] << 7) +
      (src007[69] << 7) +
      (src007[70] << 7) +
      (src007[71] << 7) +
      (src007[72] << 7) +
      (src007[73] << 7) +
      (src007[74] << 7) +
      (src007[75] << 7) +
      (src007[76] << 7) +
      (src007[77] << 7) +
      (src007[78] << 7) +
      (src007[79] << 7) +
      (src007[80] << 7) +
      (src007[81] << 7) +
      (src007[82] << 7) +
      (src007[83] << 7) +
      (src007[84] << 7) +
      (src007[85] << 7) +
      (src007[86] << 7) +
      (src007[87] << 7) +
      (src007[88] << 7) +
      (src007[89] << 7) +
      (src007[90] << 7) +
      (src007[91] << 7) +
      (src007[92] << 7) +
      (src007[93] << 7) +
      (src007[94] << 7) +
      (src007[95] << 7) +
      (src007[96] << 7) +
      (src007[97] << 7) +
      (src007[98] << 7) +
      (src007[99] << 7) +
      (src007[100] << 7) +
      (src007[101] << 7) +
      (src007[102] << 7) +
      (src007[103] << 7) +
      (src007[104] << 7) +
      (src007[105] << 7) +
      (src007[106] << 7) +
      (src007[107] << 7) +
      (src007[108] << 7) +
      (src007[109] << 7) +
      (src007[110] << 7) +
      (src007[111] << 7) +
      (src007[112] << 7) +
      (src007[113] << 7) +
      (src007[114] << 7) +
      (src007[115] << 7) +
      (src007[116] << 7) +
      (src007[117] << 7) +
      (src007[118] << 7) +
      (src007[119] << 7) +
      (src007[120] << 7) +
      (src007[121] << 7) +
      (src007[122] << 7) +
      (src007[123] << 7) +
      (src007[124] << 7) +
      (src007[125] << 7) +
      (src007[126] << 7) +
      (src007[127] << 7) +
      (src008[0] << 8) +
      (src008[1] << 8) +
      (src008[2] << 8) +
      (src008[3] << 8) +
      (src008[4] << 8) +
      (src008[5] << 8) +
      (src008[6] << 8) +
      (src008[7] << 8) +
      (src008[8] << 8) +
      (src008[9] << 8) +
      (src008[10] << 8) +
      (src008[11] << 8) +
      (src008[12] << 8) +
      (src008[13] << 8) +
      (src008[14] << 8) +
      (src008[15] << 8) +
      (src008[16] << 8) +
      (src008[17] << 8) +
      (src008[18] << 8) +
      (src008[19] << 8) +
      (src008[20] << 8) +
      (src008[21] << 8) +
      (src008[22] << 8) +
      (src008[23] << 8) +
      (src008[24] << 8) +
      (src008[25] << 8) +
      (src008[26] << 8) +
      (src008[27] << 8) +
      (src008[28] << 8) +
      (src008[29] << 8) +
      (src008[30] << 8) +
      (src008[31] << 8) +
      (src008[32] << 8) +
      (src008[33] << 8) +
      (src008[34] << 8) +
      (src008[35] << 8) +
      (src008[36] << 8) +
      (src008[37] << 8) +
      (src008[38] << 8) +
      (src008[39] << 8) +
      (src008[40] << 8) +
      (src008[41] << 8) +
      (src008[42] << 8) +
      (src008[43] << 8) +
      (src008[44] << 8) +
      (src008[45] << 8) +
      (src008[46] << 8) +
      (src008[47] << 8) +
      (src008[48] << 8) +
      (src008[49] << 8) +
      (src008[50] << 8) +
      (src008[51] << 8) +
      (src008[52] << 8) +
      (src008[53] << 8) +
      (src008[54] << 8) +
      (src008[55] << 8) +
      (src008[56] << 8) +
      (src008[57] << 8) +
      (src008[58] << 8) +
      (src008[59] << 8) +
      (src008[60] << 8) +
      (src008[61] << 8) +
      (src008[62] << 8) +
      (src008[63] << 8) +
      (src008[64] << 8) +
      (src008[65] << 8) +
      (src008[66] << 8) +
      (src008[67] << 8) +
      (src008[68] << 8) +
      (src008[69] << 8) +
      (src008[70] << 8) +
      (src008[71] << 8) +
      (src008[72] << 8) +
      (src008[73] << 8) +
      (src008[74] << 8) +
      (src008[75] << 8) +
      (src008[76] << 8) +
      (src008[77] << 8) +
      (src008[78] << 8) +
      (src008[79] << 8) +
      (src008[80] << 8) +
      (src008[81] << 8) +
      (src008[82] << 8) +
      (src008[83] << 8) +
      (src008[84] << 8) +
      (src008[85] << 8) +
      (src008[86] << 8) +
      (src008[87] << 8) +
      (src008[88] << 8) +
      (src008[89] << 8) +
      (src008[90] << 8) +
      (src008[91] << 8) +
      (src008[92] << 8) +
      (src008[93] << 8) +
      (src008[94] << 8) +
      (src008[95] << 8) +
      (src008[96] << 8) +
      (src008[97] << 8) +
      (src008[98] << 8) +
      (src008[99] << 8) +
      (src008[100] << 8) +
      (src008[101] << 8) +
      (src008[102] << 8) +
      (src008[103] << 8) +
      (src008[104] << 8) +
      (src008[105] << 8) +
      (src008[106] << 8) +
      (src008[107] << 8) +
      (src008[108] << 8) +
      (src008[109] << 8) +
      (src008[110] << 8) +
      (src008[111] << 8) +
      (src008[112] << 8) +
      (src008[113] << 8) +
      (src008[114] << 8) +
      (src008[115] << 8) +
      (src008[116] << 8) +
      (src008[117] << 8) +
      (src008[118] << 8) +
      (src008[119] << 8) +
      (src008[120] << 8) +
      (src008[121] << 8) +
      (src008[122] << 8) +
      (src008[123] << 8) +
      (src008[124] << 8) +
      (src008[125] << 8) +
      (src008[126] << 8) +
      (src008[127] << 8) +
      (src009[0] << 9) +
      (src009[1] << 9) +
      (src009[2] << 9) +
      (src009[3] << 9) +
      (src009[4] << 9) +
      (src009[5] << 9) +
      (src009[6] << 9) +
      (src009[7] << 9) +
      (src009[8] << 9) +
      (src009[9] << 9) +
      (src009[10] << 9) +
      (src009[11] << 9) +
      (src009[12] << 9) +
      (src009[13] << 9) +
      (src009[14] << 9) +
      (src009[15] << 9) +
      (src009[16] << 9) +
      (src009[17] << 9) +
      (src009[18] << 9) +
      (src009[19] << 9) +
      (src009[20] << 9) +
      (src009[21] << 9) +
      (src009[22] << 9) +
      (src009[23] << 9) +
      (src009[24] << 9) +
      (src009[25] << 9) +
      (src009[26] << 9) +
      (src009[27] << 9) +
      (src009[28] << 9) +
      (src009[29] << 9) +
      (src009[30] << 9) +
      (src009[31] << 9) +
      (src009[32] << 9) +
      (src009[33] << 9) +
      (src009[34] << 9) +
      (src009[35] << 9) +
      (src009[36] << 9) +
      (src009[37] << 9) +
      (src009[38] << 9) +
      (src009[39] << 9) +
      (src009[40] << 9) +
      (src009[41] << 9) +
      (src009[42] << 9) +
      (src009[43] << 9) +
      (src009[44] << 9) +
      (src009[45] << 9) +
      (src009[46] << 9) +
      (src009[47] << 9) +
      (src009[48] << 9) +
      (src009[49] << 9) +
      (src009[50] << 9) +
      (src009[51] << 9) +
      (src009[52] << 9) +
      (src009[53] << 9) +
      (src009[54] << 9) +
      (src009[55] << 9) +
      (src009[56] << 9) +
      (src009[57] << 9) +
      (src009[58] << 9) +
      (src009[59] << 9) +
      (src009[60] << 9) +
      (src009[61] << 9) +
      (src009[62] << 9) +
      (src009[63] << 9) +
      (src009[64] << 9) +
      (src009[65] << 9) +
      (src009[66] << 9) +
      (src009[67] << 9) +
      (src009[68] << 9) +
      (src009[69] << 9) +
      (src009[70] << 9) +
      (src009[71] << 9) +
      (src009[72] << 9) +
      (src009[73] << 9) +
      (src009[74] << 9) +
      (src009[75] << 9) +
      (src009[76] << 9) +
      (src009[77] << 9) +
      (src009[78] << 9) +
      (src009[79] << 9) +
      (src009[80] << 9) +
      (src009[81] << 9) +
      (src009[82] << 9) +
      (src009[83] << 9) +
      (src009[84] << 9) +
      (src009[85] << 9) +
      (src009[86] << 9) +
      (src009[87] << 9) +
      (src009[88] << 9) +
      (src009[89] << 9) +
      (src009[90] << 9) +
      (src009[91] << 9) +
      (src009[92] << 9) +
      (src009[93] << 9) +
      (src009[94] << 9) +
      (src009[95] << 9) +
      (src009[96] << 9) +
      (src009[97] << 9) +
      (src009[98] << 9) +
      (src009[99] << 9) +
      (src009[100] << 9) +
      (src009[101] << 9) +
      (src009[102] << 9) +
      (src009[103] << 9) +
      (src009[104] << 9) +
      (src009[105] << 9) +
      (src009[106] << 9) +
      (src009[107] << 9) +
      (src009[108] << 9) +
      (src009[109] << 9) +
      (src009[110] << 9) +
      (src009[111] << 9) +
      (src009[112] << 9) +
      (src009[113] << 9) +
      (src009[114] << 9) +
      (src009[115] << 9) +
      (src009[116] << 9) +
      (src009[117] << 9) +
      (src009[118] << 9) +
      (src009[119] << 9) +
      (src009[120] << 9) +
      (src009[121] << 9) +
      (src009[122] << 9) +
      (src009[123] << 9) +
      (src009[124] << 9) +
      (src009[125] << 9) +
      (src009[126] << 9) +
      (src009[127] << 9) +
      (src010[0] << 10) +
      (src010[1] << 10) +
      (src010[2] << 10) +
      (src010[3] << 10) +
      (src010[4] << 10) +
      (src010[5] << 10) +
      (src010[6] << 10) +
      (src010[7] << 10) +
      (src010[8] << 10) +
      (src010[9] << 10) +
      (src010[10] << 10) +
      (src010[11] << 10) +
      (src010[12] << 10) +
      (src010[13] << 10) +
      (src010[14] << 10) +
      (src010[15] << 10) +
      (src010[16] << 10) +
      (src010[17] << 10) +
      (src010[18] << 10) +
      (src010[19] << 10) +
      (src010[20] << 10) +
      (src010[21] << 10) +
      (src010[22] << 10) +
      (src010[23] << 10) +
      (src010[24] << 10) +
      (src010[25] << 10) +
      (src010[26] << 10) +
      (src010[27] << 10) +
      (src010[28] << 10) +
      (src010[29] << 10) +
      (src010[30] << 10) +
      (src010[31] << 10) +
      (src010[32] << 10) +
      (src010[33] << 10) +
      (src010[34] << 10) +
      (src010[35] << 10) +
      (src010[36] << 10) +
      (src010[37] << 10) +
      (src010[38] << 10) +
      (src010[39] << 10) +
      (src010[40] << 10) +
      (src010[41] << 10) +
      (src010[42] << 10) +
      (src010[43] << 10) +
      (src010[44] << 10) +
      (src010[45] << 10) +
      (src010[46] << 10) +
      (src010[47] << 10) +
      (src010[48] << 10) +
      (src010[49] << 10) +
      (src010[50] << 10) +
      (src010[51] << 10) +
      (src010[52] << 10) +
      (src010[53] << 10) +
      (src010[54] << 10) +
      (src010[55] << 10) +
      (src010[56] << 10) +
      (src010[57] << 10) +
      (src010[58] << 10) +
      (src010[59] << 10) +
      (src010[60] << 10) +
      (src010[61] << 10) +
      (src010[62] << 10) +
      (src010[63] << 10) +
      (src010[64] << 10) +
      (src010[65] << 10) +
      (src010[66] << 10) +
      (src010[67] << 10) +
      (src010[68] << 10) +
      (src010[69] << 10) +
      (src010[70] << 10) +
      (src010[71] << 10) +
      (src010[72] << 10) +
      (src010[73] << 10) +
      (src010[74] << 10) +
      (src010[75] << 10) +
      (src010[76] << 10) +
      (src010[77] << 10) +
      (src010[78] << 10) +
      (src010[79] << 10) +
      (src010[80] << 10) +
      (src010[81] << 10) +
      (src010[82] << 10) +
      (src010[83] << 10) +
      (src010[84] << 10) +
      (src010[85] << 10) +
      (src010[86] << 10) +
      (src010[87] << 10) +
      (src010[88] << 10) +
      (src010[89] << 10) +
      (src010[90] << 10) +
      (src010[91] << 10) +
      (src010[92] << 10) +
      (src010[93] << 10) +
      (src010[94] << 10) +
      (src010[95] << 10) +
      (src010[96] << 10) +
      (src010[97] << 10) +
      (src010[98] << 10) +
      (src010[99] << 10) +
      (src010[100] << 10) +
      (src010[101] << 10) +
      (src010[102] << 10) +
      (src010[103] << 10) +
      (src010[104] << 10) +
      (src010[105] << 10) +
      (src010[106] << 10) +
      (src010[107] << 10) +
      (src010[108] << 10) +
      (src010[109] << 10) +
      (src010[110] << 10) +
      (src010[111] << 10) +
      (src010[112] << 10) +
      (src010[113] << 10) +
      (src010[114] << 10) +
      (src010[115] << 10) +
      (src010[116] << 10) +
      (src010[117] << 10) +
      (src010[118] << 10) +
      (src010[119] << 10) +
      (src010[120] << 10) +
      (src010[121] << 10) +
      (src010[122] << 10) +
      (src010[123] << 10) +
      (src010[124] << 10) +
      (src010[125] << 10) +
      (src010[126] << 10) +
      (src010[127] << 10) +
      (src011[0] << 11) +
      (src011[1] << 11) +
      (src011[2] << 11) +
      (src011[3] << 11) +
      (src011[4] << 11) +
      (src011[5] << 11) +
      (src011[6] << 11) +
      (src011[7] << 11) +
      (src011[8] << 11) +
      (src011[9] << 11) +
      (src011[10] << 11) +
      (src011[11] << 11) +
      (src011[12] << 11) +
      (src011[13] << 11) +
      (src011[14] << 11) +
      (src011[15] << 11) +
      (src011[16] << 11) +
      (src011[17] << 11) +
      (src011[18] << 11) +
      (src011[19] << 11) +
      (src011[20] << 11) +
      (src011[21] << 11) +
      (src011[22] << 11) +
      (src011[23] << 11) +
      (src011[24] << 11) +
      (src011[25] << 11) +
      (src011[26] << 11) +
      (src011[27] << 11) +
      (src011[28] << 11) +
      (src011[29] << 11) +
      (src011[30] << 11) +
      (src011[31] << 11) +
      (src011[32] << 11) +
      (src011[33] << 11) +
      (src011[34] << 11) +
      (src011[35] << 11) +
      (src011[36] << 11) +
      (src011[37] << 11) +
      (src011[38] << 11) +
      (src011[39] << 11) +
      (src011[40] << 11) +
      (src011[41] << 11) +
      (src011[42] << 11) +
      (src011[43] << 11) +
      (src011[44] << 11) +
      (src011[45] << 11) +
      (src011[46] << 11) +
      (src011[47] << 11) +
      (src011[48] << 11) +
      (src011[49] << 11) +
      (src011[50] << 11) +
      (src011[51] << 11) +
      (src011[52] << 11) +
      (src011[53] << 11) +
      (src011[54] << 11) +
      (src011[55] << 11) +
      (src011[56] << 11) +
      (src011[57] << 11) +
      (src011[58] << 11) +
      (src011[59] << 11) +
      (src011[60] << 11) +
      (src011[61] << 11) +
      (src011[62] << 11) +
      (src011[63] << 11) +
      (src011[64] << 11) +
      (src011[65] << 11) +
      (src011[66] << 11) +
      (src011[67] << 11) +
      (src011[68] << 11) +
      (src011[69] << 11) +
      (src011[70] << 11) +
      (src011[71] << 11) +
      (src011[72] << 11) +
      (src011[73] << 11) +
      (src011[74] << 11) +
      (src011[75] << 11) +
      (src011[76] << 11) +
      (src011[77] << 11) +
      (src011[78] << 11) +
      (src011[79] << 11) +
      (src011[80] << 11) +
      (src011[81] << 11) +
      (src011[82] << 11) +
      (src011[83] << 11) +
      (src011[84] << 11) +
      (src011[85] << 11) +
      (src011[86] << 11) +
      (src011[87] << 11) +
      (src011[88] << 11) +
      (src011[89] << 11) +
      (src011[90] << 11) +
      (src011[91] << 11) +
      (src011[92] << 11) +
      (src011[93] << 11) +
      (src011[94] << 11) +
      (src011[95] << 11) +
      (src011[96] << 11) +
      (src011[97] << 11) +
      (src011[98] << 11) +
      (src011[99] << 11) +
      (src011[100] << 11) +
      (src011[101] << 11) +
      (src011[102] << 11) +
      (src011[103] << 11) +
      (src011[104] << 11) +
      (src011[105] << 11) +
      (src011[106] << 11) +
      (src011[107] << 11) +
      (src011[108] << 11) +
      (src011[109] << 11) +
      (src011[110] << 11) +
      (src011[111] << 11) +
      (src011[112] << 11) +
      (src011[113] << 11) +
      (src011[114] << 11) +
      (src011[115] << 11) +
      (src011[116] << 11) +
      (src011[117] << 11) +
      (src011[118] << 11) +
      (src011[119] << 11) +
      (src011[120] << 11) +
      (src011[121] << 11) +
      (src011[122] << 11) +
      (src011[123] << 11) +
      (src011[124] << 11) +
      (src011[125] << 11) +
      (src011[126] << 11) +
      (src011[127] << 11) +
      (src012[0] << 12) +
      (src012[1] << 12) +
      (src012[2] << 12) +
      (src012[3] << 12) +
      (src012[4] << 12) +
      (src012[5] << 12) +
      (src012[6] << 12) +
      (src012[7] << 12) +
      (src012[8] << 12) +
      (src012[9] << 12) +
      (src012[10] << 12) +
      (src012[11] << 12) +
      (src012[12] << 12) +
      (src012[13] << 12) +
      (src012[14] << 12) +
      (src012[15] << 12) +
      (src012[16] << 12) +
      (src012[17] << 12) +
      (src012[18] << 12) +
      (src012[19] << 12) +
      (src012[20] << 12) +
      (src012[21] << 12) +
      (src012[22] << 12) +
      (src012[23] << 12) +
      (src012[24] << 12) +
      (src012[25] << 12) +
      (src012[26] << 12) +
      (src012[27] << 12) +
      (src012[28] << 12) +
      (src012[29] << 12) +
      (src012[30] << 12) +
      (src012[31] << 12) +
      (src012[32] << 12) +
      (src012[33] << 12) +
      (src012[34] << 12) +
      (src012[35] << 12) +
      (src012[36] << 12) +
      (src012[37] << 12) +
      (src012[38] << 12) +
      (src012[39] << 12) +
      (src012[40] << 12) +
      (src012[41] << 12) +
      (src012[42] << 12) +
      (src012[43] << 12) +
      (src012[44] << 12) +
      (src012[45] << 12) +
      (src012[46] << 12) +
      (src012[47] << 12) +
      (src012[48] << 12) +
      (src012[49] << 12) +
      (src012[50] << 12) +
      (src012[51] << 12) +
      (src012[52] << 12) +
      (src012[53] << 12) +
      (src012[54] << 12) +
      (src012[55] << 12) +
      (src012[56] << 12) +
      (src012[57] << 12) +
      (src012[58] << 12) +
      (src012[59] << 12) +
      (src012[60] << 12) +
      (src012[61] << 12) +
      (src012[62] << 12) +
      (src012[63] << 12) +
      (src012[64] << 12) +
      (src012[65] << 12) +
      (src012[66] << 12) +
      (src012[67] << 12) +
      (src012[68] << 12) +
      (src012[69] << 12) +
      (src012[70] << 12) +
      (src012[71] << 12) +
      (src012[72] << 12) +
      (src012[73] << 12) +
      (src012[74] << 12) +
      (src012[75] << 12) +
      (src012[76] << 12) +
      (src012[77] << 12) +
      (src012[78] << 12) +
      (src012[79] << 12) +
      (src012[80] << 12) +
      (src012[81] << 12) +
      (src012[82] << 12) +
      (src012[83] << 12) +
      (src012[84] << 12) +
      (src012[85] << 12) +
      (src012[86] << 12) +
      (src012[87] << 12) +
      (src012[88] << 12) +
      (src012[89] << 12) +
      (src012[90] << 12) +
      (src012[91] << 12) +
      (src012[92] << 12) +
      (src012[93] << 12) +
      (src012[94] << 12) +
      (src012[95] << 12) +
      (src012[96] << 12) +
      (src012[97] << 12) +
      (src012[98] << 12) +
      (src012[99] << 12) +
      (src012[100] << 12) +
      (src012[101] << 12) +
      (src012[102] << 12) +
      (src012[103] << 12) +
      (src012[104] << 12) +
      (src012[105] << 12) +
      (src012[106] << 12) +
      (src012[107] << 12) +
      (src012[108] << 12) +
      (src012[109] << 12) +
      (src012[110] << 12) +
      (src012[111] << 12) +
      (src012[112] << 12) +
      (src012[113] << 12) +
      (src012[114] << 12) +
      (src012[115] << 12) +
      (src012[116] << 12) +
      (src012[117] << 12) +
      (src012[118] << 12) +
      (src012[119] << 12) +
      (src012[120] << 12) +
      (src012[121] << 12) +
      (src012[122] << 12) +
      (src012[123] << 12) +
      (src012[124] << 12) +
      (src012[125] << 12) +
      (src012[126] << 12) +
      (src012[127] << 12) +
      (src013[0] << 13) +
      (src013[1] << 13) +
      (src013[2] << 13) +
      (src013[3] << 13) +
      (src013[4] << 13) +
      (src013[5] << 13) +
      (src013[6] << 13) +
      (src013[7] << 13) +
      (src013[8] << 13) +
      (src013[9] << 13) +
      (src013[10] << 13) +
      (src013[11] << 13) +
      (src013[12] << 13) +
      (src013[13] << 13) +
      (src013[14] << 13) +
      (src013[15] << 13) +
      (src013[16] << 13) +
      (src013[17] << 13) +
      (src013[18] << 13) +
      (src013[19] << 13) +
      (src013[20] << 13) +
      (src013[21] << 13) +
      (src013[22] << 13) +
      (src013[23] << 13) +
      (src013[24] << 13) +
      (src013[25] << 13) +
      (src013[26] << 13) +
      (src013[27] << 13) +
      (src013[28] << 13) +
      (src013[29] << 13) +
      (src013[30] << 13) +
      (src013[31] << 13) +
      (src013[32] << 13) +
      (src013[33] << 13) +
      (src013[34] << 13) +
      (src013[35] << 13) +
      (src013[36] << 13) +
      (src013[37] << 13) +
      (src013[38] << 13) +
      (src013[39] << 13) +
      (src013[40] << 13) +
      (src013[41] << 13) +
      (src013[42] << 13) +
      (src013[43] << 13) +
      (src013[44] << 13) +
      (src013[45] << 13) +
      (src013[46] << 13) +
      (src013[47] << 13) +
      (src013[48] << 13) +
      (src013[49] << 13) +
      (src013[50] << 13) +
      (src013[51] << 13) +
      (src013[52] << 13) +
      (src013[53] << 13) +
      (src013[54] << 13) +
      (src013[55] << 13) +
      (src013[56] << 13) +
      (src013[57] << 13) +
      (src013[58] << 13) +
      (src013[59] << 13) +
      (src013[60] << 13) +
      (src013[61] << 13) +
      (src013[62] << 13) +
      (src013[63] << 13) +
      (src013[64] << 13) +
      (src013[65] << 13) +
      (src013[66] << 13) +
      (src013[67] << 13) +
      (src013[68] << 13) +
      (src013[69] << 13) +
      (src013[70] << 13) +
      (src013[71] << 13) +
      (src013[72] << 13) +
      (src013[73] << 13) +
      (src013[74] << 13) +
      (src013[75] << 13) +
      (src013[76] << 13) +
      (src013[77] << 13) +
      (src013[78] << 13) +
      (src013[79] << 13) +
      (src013[80] << 13) +
      (src013[81] << 13) +
      (src013[82] << 13) +
      (src013[83] << 13) +
      (src013[84] << 13) +
      (src013[85] << 13) +
      (src013[86] << 13) +
      (src013[87] << 13) +
      (src013[88] << 13) +
      (src013[89] << 13) +
      (src013[90] << 13) +
      (src013[91] << 13) +
      (src013[92] << 13) +
      (src013[93] << 13) +
      (src013[94] << 13) +
      (src013[95] << 13) +
      (src013[96] << 13) +
      (src013[97] << 13) +
      (src013[98] << 13) +
      (src013[99] << 13) +
      (src013[100] << 13) +
      (src013[101] << 13) +
      (src013[102] << 13) +
      (src013[103] << 13) +
      (src013[104] << 13) +
      (src013[105] << 13) +
      (src013[106] << 13) +
      (src013[107] << 13) +
      (src013[108] << 13) +
      (src013[109] << 13) +
      (src013[110] << 13) +
      (src013[111] << 13) +
      (src013[112] << 13) +
      (src013[113] << 13) +
      (src013[114] << 13) +
      (src013[115] << 13) +
      (src013[116] << 13) +
      (src013[117] << 13) +
      (src013[118] << 13) +
      (src013[119] << 13) +
      (src013[120] << 13) +
      (src013[121] << 13) +
      (src013[122] << 13) +
      (src013[123] << 13) +
      (src013[124] << 13) +
      (src013[125] << 13) +
      (src013[126] << 13) +
      (src013[127] << 13) +
      (src014[0] << 14) +
      (src014[1] << 14) +
      (src014[2] << 14) +
      (src014[3] << 14) +
      (src014[4] << 14) +
      (src014[5] << 14) +
      (src014[6] << 14) +
      (src014[7] << 14) +
      (src014[8] << 14) +
      (src014[9] << 14) +
      (src014[10] << 14) +
      (src014[11] << 14) +
      (src014[12] << 14) +
      (src014[13] << 14) +
      (src014[14] << 14) +
      (src014[15] << 14) +
      (src014[16] << 14) +
      (src014[17] << 14) +
      (src014[18] << 14) +
      (src014[19] << 14) +
      (src014[20] << 14) +
      (src014[21] << 14) +
      (src014[22] << 14) +
      (src014[23] << 14) +
      (src014[24] << 14) +
      (src014[25] << 14) +
      (src014[26] << 14) +
      (src014[27] << 14) +
      (src014[28] << 14) +
      (src014[29] << 14) +
      (src014[30] << 14) +
      (src014[31] << 14) +
      (src014[32] << 14) +
      (src014[33] << 14) +
      (src014[34] << 14) +
      (src014[35] << 14) +
      (src014[36] << 14) +
      (src014[37] << 14) +
      (src014[38] << 14) +
      (src014[39] << 14) +
      (src014[40] << 14) +
      (src014[41] << 14) +
      (src014[42] << 14) +
      (src014[43] << 14) +
      (src014[44] << 14) +
      (src014[45] << 14) +
      (src014[46] << 14) +
      (src014[47] << 14) +
      (src014[48] << 14) +
      (src014[49] << 14) +
      (src014[50] << 14) +
      (src014[51] << 14) +
      (src014[52] << 14) +
      (src014[53] << 14) +
      (src014[54] << 14) +
      (src014[55] << 14) +
      (src014[56] << 14) +
      (src014[57] << 14) +
      (src014[58] << 14) +
      (src014[59] << 14) +
      (src014[60] << 14) +
      (src014[61] << 14) +
      (src014[62] << 14) +
      (src014[63] << 14) +
      (src014[64] << 14) +
      (src014[65] << 14) +
      (src014[66] << 14) +
      (src014[67] << 14) +
      (src014[68] << 14) +
      (src014[69] << 14) +
      (src014[70] << 14) +
      (src014[71] << 14) +
      (src014[72] << 14) +
      (src014[73] << 14) +
      (src014[74] << 14) +
      (src014[75] << 14) +
      (src014[76] << 14) +
      (src014[77] << 14) +
      (src014[78] << 14) +
      (src014[79] << 14) +
      (src014[80] << 14) +
      (src014[81] << 14) +
      (src014[82] << 14) +
      (src014[83] << 14) +
      (src014[84] << 14) +
      (src014[85] << 14) +
      (src014[86] << 14) +
      (src014[87] << 14) +
      (src014[88] << 14) +
      (src014[89] << 14) +
      (src014[90] << 14) +
      (src014[91] << 14) +
      (src014[92] << 14) +
      (src014[93] << 14) +
      (src014[94] << 14) +
      (src014[95] << 14) +
      (src014[96] << 14) +
      (src014[97] << 14) +
      (src014[98] << 14) +
      (src014[99] << 14) +
      (src014[100] << 14) +
      (src014[101] << 14) +
      (src014[102] << 14) +
      (src014[103] << 14) +
      (src014[104] << 14) +
      (src014[105] << 14) +
      (src014[106] << 14) +
      (src014[107] << 14) +
      (src014[108] << 14) +
      (src014[109] << 14) +
      (src014[110] << 14) +
      (src014[111] << 14) +
      (src014[112] << 14) +
      (src014[113] << 14) +
      (src014[114] << 14) +
      (src014[115] << 14) +
      (src014[116] << 14) +
      (src014[117] << 14) +
      (src014[118] << 14) +
      (src014[119] << 14) +
      (src014[120] << 14) +
      (src014[121] << 14) +
      (src014[122] << 14) +
      (src014[123] << 14) +
      (src014[124] << 14) +
      (src014[125] << 14) +
      (src014[126] << 14) +
      (src014[127] << 14) +
      (src015[0] << 15) +
      (src015[1] << 15) +
      (src015[2] << 15) +
      (src015[3] << 15) +
      (src015[4] << 15) +
      (src015[5] << 15) +
      (src015[6] << 15) +
      (src015[7] << 15) +
      (src015[8] << 15) +
      (src015[9] << 15) +
      (src015[10] << 15) +
      (src015[11] << 15) +
      (src015[12] << 15) +
      (src015[13] << 15) +
      (src015[14] << 15) +
      (src015[15] << 15) +
      (src015[16] << 15) +
      (src015[17] << 15) +
      (src015[18] << 15) +
      (src015[19] << 15) +
      (src015[20] << 15) +
      (src015[21] << 15) +
      (src015[22] << 15) +
      (src015[23] << 15) +
      (src015[24] << 15) +
      (src015[25] << 15) +
      (src015[26] << 15) +
      (src015[27] << 15) +
      (src015[28] << 15) +
      (src015[29] << 15) +
      (src015[30] << 15) +
      (src015[31] << 15) +
      (src015[32] << 15) +
      (src015[33] << 15) +
      (src015[34] << 15) +
      (src015[35] << 15) +
      (src015[36] << 15) +
      (src015[37] << 15) +
      (src015[38] << 15) +
      (src015[39] << 15) +
      (src015[40] << 15) +
      (src015[41] << 15) +
      (src015[42] << 15) +
      (src015[43] << 15) +
      (src015[44] << 15) +
      (src015[45] << 15) +
      (src015[46] << 15) +
      (src015[47] << 15) +
      (src015[48] << 15) +
      (src015[49] << 15) +
      (src015[50] << 15) +
      (src015[51] << 15) +
      (src015[52] << 15) +
      (src015[53] << 15) +
      (src015[54] << 15) +
      (src015[55] << 15) +
      (src015[56] << 15) +
      (src015[57] << 15) +
      (src015[58] << 15) +
      (src015[59] << 15) +
      (src015[60] << 15) +
      (src015[61] << 15) +
      (src015[62] << 15) +
      (src015[63] << 15) +
      (src015[64] << 15) +
      (src015[65] << 15) +
      (src015[66] << 15) +
      (src015[67] << 15) +
      (src015[68] << 15) +
      (src015[69] << 15) +
      (src015[70] << 15) +
      (src015[71] << 15) +
      (src015[72] << 15) +
      (src015[73] << 15) +
      (src015[74] << 15) +
      (src015[75] << 15) +
      (src015[76] << 15) +
      (src015[77] << 15) +
      (src015[78] << 15) +
      (src015[79] << 15) +
      (src015[80] << 15) +
      (src015[81] << 15) +
      (src015[82] << 15) +
      (src015[83] << 15) +
      (src015[84] << 15) +
      (src015[85] << 15) +
      (src015[86] << 15) +
      (src015[87] << 15) +
      (src015[88] << 15) +
      (src015[89] << 15) +
      (src015[90] << 15) +
      (src015[91] << 15) +
      (src015[92] << 15) +
      (src015[93] << 15) +
      (src015[94] << 15) +
      (src015[95] << 15) +
      (src015[96] << 15) +
      (src015[97] << 15) +
      (src015[98] << 15) +
      (src015[99] << 15) +
      (src015[100] << 15) +
      (src015[101] << 15) +
      (src015[102] << 15) +
      (src015[103] << 15) +
      (src015[104] << 15) +
      (src015[105] << 15) +
      (src015[106] << 15) +
      (src015[107] << 15) +
      (src015[108] << 15) +
      (src015[109] << 15) +
      (src015[110] << 15) +
      (src015[111] << 15) +
      (src015[112] << 15) +
      (src015[113] << 15) +
      (src015[114] << 15) +
      (src015[115] << 15) +
      (src015[116] << 15) +
      (src015[117] << 15) +
      (src015[118] << 15) +
      (src015[119] << 15) +
      (src015[120] << 15) +
      (src015[121] << 15) +
      (src015[122] << 15) +
      (src015[123] << 15) +
      (src015[124] << 15) +
      (src015[125] << 15) +
      (src015[126] << 15) +
      (src015[127] << 15) +
      (src016[0] << 16) +
      (src016[1] << 16) +
      (src016[2] << 16) +
      (src016[3] << 16) +
      (src016[4] << 16) +
      (src016[5] << 16) +
      (src016[6] << 16) +
      (src016[7] << 16) +
      (src016[8] << 16) +
      (src016[9] << 16) +
      (src016[10] << 16) +
      (src016[11] << 16) +
      (src016[12] << 16) +
      (src016[13] << 16) +
      (src016[14] << 16) +
      (src016[15] << 16) +
      (src016[16] << 16) +
      (src016[17] << 16) +
      (src016[18] << 16) +
      (src016[19] << 16) +
      (src016[20] << 16) +
      (src016[21] << 16) +
      (src016[22] << 16) +
      (src016[23] << 16) +
      (src016[24] << 16) +
      (src016[25] << 16) +
      (src016[26] << 16) +
      (src016[27] << 16) +
      (src016[28] << 16) +
      (src016[29] << 16) +
      (src016[30] << 16) +
      (src016[31] << 16) +
      (src016[32] << 16) +
      (src016[33] << 16) +
      (src016[34] << 16) +
      (src016[35] << 16) +
      (src016[36] << 16) +
      (src016[37] << 16) +
      (src016[38] << 16) +
      (src016[39] << 16) +
      (src016[40] << 16) +
      (src016[41] << 16) +
      (src016[42] << 16) +
      (src016[43] << 16) +
      (src016[44] << 16) +
      (src016[45] << 16) +
      (src016[46] << 16) +
      (src016[47] << 16) +
      (src016[48] << 16) +
      (src016[49] << 16) +
      (src016[50] << 16) +
      (src016[51] << 16) +
      (src016[52] << 16) +
      (src016[53] << 16) +
      (src016[54] << 16) +
      (src016[55] << 16) +
      (src016[56] << 16) +
      (src016[57] << 16) +
      (src016[58] << 16) +
      (src016[59] << 16) +
      (src016[60] << 16) +
      (src016[61] << 16) +
      (src016[62] << 16) +
      (src016[63] << 16) +
      (src016[64] << 16) +
      (src016[65] << 16) +
      (src016[66] << 16) +
      (src016[67] << 16) +
      (src016[68] << 16) +
      (src016[69] << 16) +
      (src016[70] << 16) +
      (src016[71] << 16) +
      (src016[72] << 16) +
      (src016[73] << 16) +
      (src016[74] << 16) +
      (src016[75] << 16) +
      (src016[76] << 16) +
      (src016[77] << 16) +
      (src016[78] << 16) +
      (src016[79] << 16) +
      (src016[80] << 16) +
      (src016[81] << 16) +
      (src016[82] << 16) +
      (src016[83] << 16) +
      (src016[84] << 16) +
      (src016[85] << 16) +
      (src016[86] << 16) +
      (src016[87] << 16) +
      (src016[88] << 16) +
      (src016[89] << 16) +
      (src016[90] << 16) +
      (src016[91] << 16) +
      (src016[92] << 16) +
      (src016[93] << 16) +
      (src016[94] << 16) +
      (src016[95] << 16) +
      (src016[96] << 16) +
      (src016[97] << 16) +
      (src016[98] << 16) +
      (src016[99] << 16) +
      (src016[100] << 16) +
      (src016[101] << 16) +
      (src016[102] << 16) +
      (src016[103] << 16) +
      (src016[104] << 16) +
      (src016[105] << 16) +
      (src016[106] << 16) +
      (src016[107] << 16) +
      (src016[108] << 16) +
      (src016[109] << 16) +
      (src016[110] << 16) +
      (src016[111] << 16) +
      (src016[112] << 16) +
      (src016[113] << 16) +
      (src016[114] << 16) +
      (src016[115] << 16) +
      (src016[116] << 16) +
      (src016[117] << 16) +
      (src016[118] << 16) +
      (src016[119] << 16) +
      (src016[120] << 16) +
      (src016[121] << 16) +
      (src016[122] << 16) +
      (src016[123] << 16) +
      (src016[124] << 16) +
      (src016[125] << 16) +
      (src016[126] << 16) +
      (src016[127] << 16) +
      (src017[0] << 17) +
      (src017[1] << 17) +
      (src017[2] << 17) +
      (src017[3] << 17) +
      (src017[4] << 17) +
      (src017[5] << 17) +
      (src017[6] << 17) +
      (src017[7] << 17) +
      (src017[8] << 17) +
      (src017[9] << 17) +
      (src017[10] << 17) +
      (src017[11] << 17) +
      (src017[12] << 17) +
      (src017[13] << 17) +
      (src017[14] << 17) +
      (src017[15] << 17) +
      (src017[16] << 17) +
      (src017[17] << 17) +
      (src017[18] << 17) +
      (src017[19] << 17) +
      (src017[20] << 17) +
      (src017[21] << 17) +
      (src017[22] << 17) +
      (src017[23] << 17) +
      (src017[24] << 17) +
      (src017[25] << 17) +
      (src017[26] << 17) +
      (src017[27] << 17) +
      (src017[28] << 17) +
      (src017[29] << 17) +
      (src017[30] << 17) +
      (src017[31] << 17) +
      (src017[32] << 17) +
      (src017[33] << 17) +
      (src017[34] << 17) +
      (src017[35] << 17) +
      (src017[36] << 17) +
      (src017[37] << 17) +
      (src017[38] << 17) +
      (src017[39] << 17) +
      (src017[40] << 17) +
      (src017[41] << 17) +
      (src017[42] << 17) +
      (src017[43] << 17) +
      (src017[44] << 17) +
      (src017[45] << 17) +
      (src017[46] << 17) +
      (src017[47] << 17) +
      (src017[48] << 17) +
      (src017[49] << 17) +
      (src017[50] << 17) +
      (src017[51] << 17) +
      (src017[52] << 17) +
      (src017[53] << 17) +
      (src017[54] << 17) +
      (src017[55] << 17) +
      (src017[56] << 17) +
      (src017[57] << 17) +
      (src017[58] << 17) +
      (src017[59] << 17) +
      (src017[60] << 17) +
      (src017[61] << 17) +
      (src017[62] << 17) +
      (src017[63] << 17) +
      (src017[64] << 17) +
      (src017[65] << 17) +
      (src017[66] << 17) +
      (src017[67] << 17) +
      (src017[68] << 17) +
      (src017[69] << 17) +
      (src017[70] << 17) +
      (src017[71] << 17) +
      (src017[72] << 17) +
      (src017[73] << 17) +
      (src017[74] << 17) +
      (src017[75] << 17) +
      (src017[76] << 17) +
      (src017[77] << 17) +
      (src017[78] << 17) +
      (src017[79] << 17) +
      (src017[80] << 17) +
      (src017[81] << 17) +
      (src017[82] << 17) +
      (src017[83] << 17) +
      (src017[84] << 17) +
      (src017[85] << 17) +
      (src017[86] << 17) +
      (src017[87] << 17) +
      (src017[88] << 17) +
      (src017[89] << 17) +
      (src017[90] << 17) +
      (src017[91] << 17) +
      (src017[92] << 17) +
      (src017[93] << 17) +
      (src017[94] << 17) +
      (src017[95] << 17) +
      (src017[96] << 17) +
      (src017[97] << 17) +
      (src017[98] << 17) +
      (src017[99] << 17) +
      (src017[100] << 17) +
      (src017[101] << 17) +
      (src017[102] << 17) +
      (src017[103] << 17) +
      (src017[104] << 17) +
      (src017[105] << 17) +
      (src017[106] << 17) +
      (src017[107] << 17) +
      (src017[108] << 17) +
      (src017[109] << 17) +
      (src017[110] << 17) +
      (src017[111] << 17) +
      (src017[112] << 17) +
      (src017[113] << 17) +
      (src017[114] << 17) +
      (src017[115] << 17) +
      (src017[116] << 17) +
      (src017[117] << 17) +
      (src017[118] << 17) +
      (src017[119] << 17) +
      (src017[120] << 17) +
      (src017[121] << 17) +
      (src017[122] << 17) +
      (src017[123] << 17) +
      (src017[124] << 17) +
      (src017[125] << 17) +
      (src017[126] << 17) +
      (src017[127] << 17) +
      (src018[0] << 18) +
      (src018[1] << 18) +
      (src018[2] << 18) +
      (src018[3] << 18) +
      (src018[4] << 18) +
      (src018[5] << 18) +
      (src018[6] << 18) +
      (src018[7] << 18) +
      (src018[8] << 18) +
      (src018[9] << 18) +
      (src018[10] << 18) +
      (src018[11] << 18) +
      (src018[12] << 18) +
      (src018[13] << 18) +
      (src018[14] << 18) +
      (src018[15] << 18) +
      (src018[16] << 18) +
      (src018[17] << 18) +
      (src018[18] << 18) +
      (src018[19] << 18) +
      (src018[20] << 18) +
      (src018[21] << 18) +
      (src018[22] << 18) +
      (src018[23] << 18) +
      (src018[24] << 18) +
      (src018[25] << 18) +
      (src018[26] << 18) +
      (src018[27] << 18) +
      (src018[28] << 18) +
      (src018[29] << 18) +
      (src018[30] << 18) +
      (src018[31] << 18) +
      (src018[32] << 18) +
      (src018[33] << 18) +
      (src018[34] << 18) +
      (src018[35] << 18) +
      (src018[36] << 18) +
      (src018[37] << 18) +
      (src018[38] << 18) +
      (src018[39] << 18) +
      (src018[40] << 18) +
      (src018[41] << 18) +
      (src018[42] << 18) +
      (src018[43] << 18) +
      (src018[44] << 18) +
      (src018[45] << 18) +
      (src018[46] << 18) +
      (src018[47] << 18) +
      (src018[48] << 18) +
      (src018[49] << 18) +
      (src018[50] << 18) +
      (src018[51] << 18) +
      (src018[52] << 18) +
      (src018[53] << 18) +
      (src018[54] << 18) +
      (src018[55] << 18) +
      (src018[56] << 18) +
      (src018[57] << 18) +
      (src018[58] << 18) +
      (src018[59] << 18) +
      (src018[60] << 18) +
      (src018[61] << 18) +
      (src018[62] << 18) +
      (src018[63] << 18) +
      (src018[64] << 18) +
      (src018[65] << 18) +
      (src018[66] << 18) +
      (src018[67] << 18) +
      (src018[68] << 18) +
      (src018[69] << 18) +
      (src018[70] << 18) +
      (src018[71] << 18) +
      (src018[72] << 18) +
      (src018[73] << 18) +
      (src018[74] << 18) +
      (src018[75] << 18) +
      (src018[76] << 18) +
      (src018[77] << 18) +
      (src018[78] << 18) +
      (src018[79] << 18) +
      (src018[80] << 18) +
      (src018[81] << 18) +
      (src018[82] << 18) +
      (src018[83] << 18) +
      (src018[84] << 18) +
      (src018[85] << 18) +
      (src018[86] << 18) +
      (src018[87] << 18) +
      (src018[88] << 18) +
      (src018[89] << 18) +
      (src018[90] << 18) +
      (src018[91] << 18) +
      (src018[92] << 18) +
      (src018[93] << 18) +
      (src018[94] << 18) +
      (src018[95] << 18) +
      (src018[96] << 18) +
      (src018[97] << 18) +
      (src018[98] << 18) +
      (src018[99] << 18) +
      (src018[100] << 18) +
      (src018[101] << 18) +
      (src018[102] << 18) +
      (src018[103] << 18) +
      (src018[104] << 18) +
      (src018[105] << 18) +
      (src018[106] << 18) +
      (src018[107] << 18) +
      (src018[108] << 18) +
      (src018[109] << 18) +
      (src018[110] << 18) +
      (src018[111] << 18) +
      (src018[112] << 18) +
      (src018[113] << 18) +
      (src018[114] << 18) +
      (src018[115] << 18) +
      (src018[116] << 18) +
      (src018[117] << 18) +
      (src018[118] << 18) +
      (src018[119] << 18) +
      (src018[120] << 18) +
      (src018[121] << 18) +
      (src018[122] << 18) +
      (src018[123] << 18) +
      (src018[124] << 18) +
      (src018[125] << 18) +
      (src018[126] << 18) +
      (src018[127] << 18) +
      (src019[0] << 19) +
      (src019[1] << 19) +
      (src019[2] << 19) +
      (src019[3] << 19) +
      (src019[4] << 19) +
      (src019[5] << 19) +
      (src019[6] << 19) +
      (src019[7] << 19) +
      (src019[8] << 19) +
      (src019[9] << 19) +
      (src019[10] << 19) +
      (src019[11] << 19) +
      (src019[12] << 19) +
      (src019[13] << 19) +
      (src019[14] << 19) +
      (src019[15] << 19) +
      (src019[16] << 19) +
      (src019[17] << 19) +
      (src019[18] << 19) +
      (src019[19] << 19) +
      (src019[20] << 19) +
      (src019[21] << 19) +
      (src019[22] << 19) +
      (src019[23] << 19) +
      (src019[24] << 19) +
      (src019[25] << 19) +
      (src019[26] << 19) +
      (src019[27] << 19) +
      (src019[28] << 19) +
      (src019[29] << 19) +
      (src019[30] << 19) +
      (src019[31] << 19) +
      (src019[32] << 19) +
      (src019[33] << 19) +
      (src019[34] << 19) +
      (src019[35] << 19) +
      (src019[36] << 19) +
      (src019[37] << 19) +
      (src019[38] << 19) +
      (src019[39] << 19) +
      (src019[40] << 19) +
      (src019[41] << 19) +
      (src019[42] << 19) +
      (src019[43] << 19) +
      (src019[44] << 19) +
      (src019[45] << 19) +
      (src019[46] << 19) +
      (src019[47] << 19) +
      (src019[48] << 19) +
      (src019[49] << 19) +
      (src019[50] << 19) +
      (src019[51] << 19) +
      (src019[52] << 19) +
      (src019[53] << 19) +
      (src019[54] << 19) +
      (src019[55] << 19) +
      (src019[56] << 19) +
      (src019[57] << 19) +
      (src019[58] << 19) +
      (src019[59] << 19) +
      (src019[60] << 19) +
      (src019[61] << 19) +
      (src019[62] << 19) +
      (src019[63] << 19) +
      (src019[64] << 19) +
      (src019[65] << 19) +
      (src019[66] << 19) +
      (src019[67] << 19) +
      (src019[68] << 19) +
      (src019[69] << 19) +
      (src019[70] << 19) +
      (src019[71] << 19) +
      (src019[72] << 19) +
      (src019[73] << 19) +
      (src019[74] << 19) +
      (src019[75] << 19) +
      (src019[76] << 19) +
      (src019[77] << 19) +
      (src019[78] << 19) +
      (src019[79] << 19) +
      (src019[80] << 19) +
      (src019[81] << 19) +
      (src019[82] << 19) +
      (src019[83] << 19) +
      (src019[84] << 19) +
      (src019[85] << 19) +
      (src019[86] << 19) +
      (src019[87] << 19) +
      (src019[88] << 19) +
      (src019[89] << 19) +
      (src019[90] << 19) +
      (src019[91] << 19) +
      (src019[92] << 19) +
      (src019[93] << 19) +
      (src019[94] << 19) +
      (src019[95] << 19) +
      (src019[96] << 19) +
      (src019[97] << 19) +
      (src019[98] << 19) +
      (src019[99] << 19) +
      (src019[100] << 19) +
      (src019[101] << 19) +
      (src019[102] << 19) +
      (src019[103] << 19) +
      (src019[104] << 19) +
      (src019[105] << 19) +
      (src019[106] << 19) +
      (src019[107] << 19) +
      (src019[108] << 19) +
      (src019[109] << 19) +
      (src019[110] << 19) +
      (src019[111] << 19) +
      (src019[112] << 19) +
      (src019[113] << 19) +
      (src019[114] << 19) +
      (src019[115] << 19) +
      (src019[116] << 19) +
      (src019[117] << 19) +
      (src019[118] << 19) +
      (src019[119] << 19) +
      (src019[120] << 19) +
      (src019[121] << 19) +
      (src019[122] << 19) +
      (src019[123] << 19) +
      (src019[124] << 19) +
      (src019[125] << 19) +
      (src019[126] << 19) +
      (src019[127] << 19) +
      (src020[0] << 20) +
      (src020[1] << 20) +
      (src020[2] << 20) +
      (src020[3] << 20) +
      (src020[4] << 20) +
      (src020[5] << 20) +
      (src020[6] << 20) +
      (src020[7] << 20) +
      (src020[8] << 20) +
      (src020[9] << 20) +
      (src020[10] << 20) +
      (src020[11] << 20) +
      (src020[12] << 20) +
      (src020[13] << 20) +
      (src020[14] << 20) +
      (src020[15] << 20) +
      (src020[16] << 20) +
      (src020[17] << 20) +
      (src020[18] << 20) +
      (src020[19] << 20) +
      (src020[20] << 20) +
      (src020[21] << 20) +
      (src020[22] << 20) +
      (src020[23] << 20) +
      (src020[24] << 20) +
      (src020[25] << 20) +
      (src020[26] << 20) +
      (src020[27] << 20) +
      (src020[28] << 20) +
      (src020[29] << 20) +
      (src020[30] << 20) +
      (src020[31] << 20) +
      (src020[32] << 20) +
      (src020[33] << 20) +
      (src020[34] << 20) +
      (src020[35] << 20) +
      (src020[36] << 20) +
      (src020[37] << 20) +
      (src020[38] << 20) +
      (src020[39] << 20) +
      (src020[40] << 20) +
      (src020[41] << 20) +
      (src020[42] << 20) +
      (src020[43] << 20) +
      (src020[44] << 20) +
      (src020[45] << 20) +
      (src020[46] << 20) +
      (src020[47] << 20) +
      (src020[48] << 20) +
      (src020[49] << 20) +
      (src020[50] << 20) +
      (src020[51] << 20) +
      (src020[52] << 20) +
      (src020[53] << 20) +
      (src020[54] << 20) +
      (src020[55] << 20) +
      (src020[56] << 20) +
      (src020[57] << 20) +
      (src020[58] << 20) +
      (src020[59] << 20) +
      (src020[60] << 20) +
      (src020[61] << 20) +
      (src020[62] << 20) +
      (src020[63] << 20) +
      (src020[64] << 20) +
      (src020[65] << 20) +
      (src020[66] << 20) +
      (src020[67] << 20) +
      (src020[68] << 20) +
      (src020[69] << 20) +
      (src020[70] << 20) +
      (src020[71] << 20) +
      (src020[72] << 20) +
      (src020[73] << 20) +
      (src020[74] << 20) +
      (src020[75] << 20) +
      (src020[76] << 20) +
      (src020[77] << 20) +
      (src020[78] << 20) +
      (src020[79] << 20) +
      (src020[80] << 20) +
      (src020[81] << 20) +
      (src020[82] << 20) +
      (src020[83] << 20) +
      (src020[84] << 20) +
      (src020[85] << 20) +
      (src020[86] << 20) +
      (src020[87] << 20) +
      (src020[88] << 20) +
      (src020[89] << 20) +
      (src020[90] << 20) +
      (src020[91] << 20) +
      (src020[92] << 20) +
      (src020[93] << 20) +
      (src020[94] << 20) +
      (src020[95] << 20) +
      (src020[96] << 20) +
      (src020[97] << 20) +
      (src020[98] << 20) +
      (src020[99] << 20) +
      (src020[100] << 20) +
      (src020[101] << 20) +
      (src020[102] << 20) +
      (src020[103] << 20) +
      (src020[104] << 20) +
      (src020[105] << 20) +
      (src020[106] << 20) +
      (src020[107] << 20) +
      (src020[108] << 20) +
      (src020[109] << 20) +
      (src020[110] << 20) +
      (src020[111] << 20) +
      (src020[112] << 20) +
      (src020[113] << 20) +
      (src020[114] << 20) +
      (src020[115] << 20) +
      (src020[116] << 20) +
      (src020[117] << 20) +
      (src020[118] << 20) +
      (src020[119] << 20) +
      (src020[120] << 20) +
      (src020[121] << 20) +
      (src020[122] << 20) +
      (src020[123] << 20) +
      (src020[124] << 20) +
      (src020[125] << 20) +
      (src020[126] << 20) +
      (src020[127] << 20) +
      (src021[0] << 21) +
      (src021[1] << 21) +
      (src021[2] << 21) +
      (src021[3] << 21) +
      (src021[4] << 21) +
      (src021[5] << 21) +
      (src021[6] << 21) +
      (src021[7] << 21) +
      (src021[8] << 21) +
      (src021[9] << 21) +
      (src021[10] << 21) +
      (src021[11] << 21) +
      (src021[12] << 21) +
      (src021[13] << 21) +
      (src021[14] << 21) +
      (src021[15] << 21) +
      (src021[16] << 21) +
      (src021[17] << 21) +
      (src021[18] << 21) +
      (src021[19] << 21) +
      (src021[20] << 21) +
      (src021[21] << 21) +
      (src021[22] << 21) +
      (src021[23] << 21) +
      (src021[24] << 21) +
      (src021[25] << 21) +
      (src021[26] << 21) +
      (src021[27] << 21) +
      (src021[28] << 21) +
      (src021[29] << 21) +
      (src021[30] << 21) +
      (src021[31] << 21) +
      (src021[32] << 21) +
      (src021[33] << 21) +
      (src021[34] << 21) +
      (src021[35] << 21) +
      (src021[36] << 21) +
      (src021[37] << 21) +
      (src021[38] << 21) +
      (src021[39] << 21) +
      (src021[40] << 21) +
      (src021[41] << 21) +
      (src021[42] << 21) +
      (src021[43] << 21) +
      (src021[44] << 21) +
      (src021[45] << 21) +
      (src021[46] << 21) +
      (src021[47] << 21) +
      (src021[48] << 21) +
      (src021[49] << 21) +
      (src021[50] << 21) +
      (src021[51] << 21) +
      (src021[52] << 21) +
      (src021[53] << 21) +
      (src021[54] << 21) +
      (src021[55] << 21) +
      (src021[56] << 21) +
      (src021[57] << 21) +
      (src021[58] << 21) +
      (src021[59] << 21) +
      (src021[60] << 21) +
      (src021[61] << 21) +
      (src021[62] << 21) +
      (src021[63] << 21) +
      (src021[64] << 21) +
      (src021[65] << 21) +
      (src021[66] << 21) +
      (src021[67] << 21) +
      (src021[68] << 21) +
      (src021[69] << 21) +
      (src021[70] << 21) +
      (src021[71] << 21) +
      (src021[72] << 21) +
      (src021[73] << 21) +
      (src021[74] << 21) +
      (src021[75] << 21) +
      (src021[76] << 21) +
      (src021[77] << 21) +
      (src021[78] << 21) +
      (src021[79] << 21) +
      (src021[80] << 21) +
      (src021[81] << 21) +
      (src021[82] << 21) +
      (src021[83] << 21) +
      (src021[84] << 21) +
      (src021[85] << 21) +
      (src021[86] << 21) +
      (src021[87] << 21) +
      (src021[88] << 21) +
      (src021[89] << 21) +
      (src021[90] << 21) +
      (src021[91] << 21) +
      (src021[92] << 21) +
      (src021[93] << 21) +
      (src021[94] << 21) +
      (src021[95] << 21) +
      (src021[96] << 21) +
      (src021[97] << 21) +
      (src021[98] << 21) +
      (src021[99] << 21) +
      (src021[100] << 21) +
      (src021[101] << 21) +
      (src021[102] << 21) +
      (src021[103] << 21) +
      (src021[104] << 21) +
      (src021[105] << 21) +
      (src021[106] << 21) +
      (src021[107] << 21) +
      (src021[108] << 21) +
      (src021[109] << 21) +
      (src021[110] << 21) +
      (src021[111] << 21) +
      (src021[112] << 21) +
      (src021[113] << 21) +
      (src021[114] << 21) +
      (src021[115] << 21) +
      (src021[116] << 21) +
      (src021[117] << 21) +
      (src021[118] << 21) +
      (src021[119] << 21) +
      (src021[120] << 21) +
      (src021[121] << 21) +
      (src021[122] << 21) +
      (src021[123] << 21) +
      (src021[124] << 21) +
      (src021[125] << 21) +
      (src021[126] << 21) +
      (src021[127] << 21) +
      (src022[0] << 22) +
      (src022[1] << 22) +
      (src022[2] << 22) +
      (src022[3] << 22) +
      (src022[4] << 22) +
      (src022[5] << 22) +
      (src022[6] << 22) +
      (src022[7] << 22) +
      (src022[8] << 22) +
      (src022[9] << 22) +
      (src022[10] << 22) +
      (src022[11] << 22) +
      (src022[12] << 22) +
      (src022[13] << 22) +
      (src022[14] << 22) +
      (src022[15] << 22) +
      (src022[16] << 22) +
      (src022[17] << 22) +
      (src022[18] << 22) +
      (src022[19] << 22) +
      (src022[20] << 22) +
      (src022[21] << 22) +
      (src022[22] << 22) +
      (src022[23] << 22) +
      (src022[24] << 22) +
      (src022[25] << 22) +
      (src022[26] << 22) +
      (src022[27] << 22) +
      (src022[28] << 22) +
      (src022[29] << 22) +
      (src022[30] << 22) +
      (src022[31] << 22) +
      (src022[32] << 22) +
      (src022[33] << 22) +
      (src022[34] << 22) +
      (src022[35] << 22) +
      (src022[36] << 22) +
      (src022[37] << 22) +
      (src022[38] << 22) +
      (src022[39] << 22) +
      (src022[40] << 22) +
      (src022[41] << 22) +
      (src022[42] << 22) +
      (src022[43] << 22) +
      (src022[44] << 22) +
      (src022[45] << 22) +
      (src022[46] << 22) +
      (src022[47] << 22) +
      (src022[48] << 22) +
      (src022[49] << 22) +
      (src022[50] << 22) +
      (src022[51] << 22) +
      (src022[52] << 22) +
      (src022[53] << 22) +
      (src022[54] << 22) +
      (src022[55] << 22) +
      (src022[56] << 22) +
      (src022[57] << 22) +
      (src022[58] << 22) +
      (src022[59] << 22) +
      (src022[60] << 22) +
      (src022[61] << 22) +
      (src022[62] << 22) +
      (src022[63] << 22) +
      (src022[64] << 22) +
      (src022[65] << 22) +
      (src022[66] << 22) +
      (src022[67] << 22) +
      (src022[68] << 22) +
      (src022[69] << 22) +
      (src022[70] << 22) +
      (src022[71] << 22) +
      (src022[72] << 22) +
      (src022[73] << 22) +
      (src022[74] << 22) +
      (src022[75] << 22) +
      (src022[76] << 22) +
      (src022[77] << 22) +
      (src022[78] << 22) +
      (src022[79] << 22) +
      (src022[80] << 22) +
      (src022[81] << 22) +
      (src022[82] << 22) +
      (src022[83] << 22) +
      (src022[84] << 22) +
      (src022[85] << 22) +
      (src022[86] << 22) +
      (src022[87] << 22) +
      (src022[88] << 22) +
      (src022[89] << 22) +
      (src022[90] << 22) +
      (src022[91] << 22) +
      (src022[92] << 22) +
      (src022[93] << 22) +
      (src022[94] << 22) +
      (src022[95] << 22) +
      (src022[96] << 22) +
      (src022[97] << 22) +
      (src022[98] << 22) +
      (src022[99] << 22) +
      (src022[100] << 22) +
      (src022[101] << 22) +
      (src022[102] << 22) +
      (src022[103] << 22) +
      (src022[104] << 22) +
      (src022[105] << 22) +
      (src022[106] << 22) +
      (src022[107] << 22) +
      (src022[108] << 22) +
      (src022[109] << 22) +
      (src022[110] << 22) +
      (src022[111] << 22) +
      (src022[112] << 22) +
      (src022[113] << 22) +
      (src022[114] << 22) +
      (src022[115] << 22) +
      (src022[116] << 22) +
      (src022[117] << 22) +
      (src022[118] << 22) +
      (src022[119] << 22) +
      (src022[120] << 22) +
      (src022[121] << 22) +
      (src022[122] << 22) +
      (src022[123] << 22) +
      (src022[124] << 22) +
      (src022[125] << 22) +
      (src022[126] << 22) +
      (src022[127] << 22) +
      (src023[0] << 23) +
      (src023[1] << 23) +
      (src023[2] << 23) +
      (src023[3] << 23) +
      (src023[4] << 23) +
      (src023[5] << 23) +
      (src023[6] << 23) +
      (src023[7] << 23) +
      (src023[8] << 23) +
      (src023[9] << 23) +
      (src023[10] << 23) +
      (src023[11] << 23) +
      (src023[12] << 23) +
      (src023[13] << 23) +
      (src023[14] << 23) +
      (src023[15] << 23) +
      (src023[16] << 23) +
      (src023[17] << 23) +
      (src023[18] << 23) +
      (src023[19] << 23) +
      (src023[20] << 23) +
      (src023[21] << 23) +
      (src023[22] << 23) +
      (src023[23] << 23) +
      (src023[24] << 23) +
      (src023[25] << 23) +
      (src023[26] << 23) +
      (src023[27] << 23) +
      (src023[28] << 23) +
      (src023[29] << 23) +
      (src023[30] << 23) +
      (src023[31] << 23) +
      (src023[32] << 23) +
      (src023[33] << 23) +
      (src023[34] << 23) +
      (src023[35] << 23) +
      (src023[36] << 23) +
      (src023[37] << 23) +
      (src023[38] << 23) +
      (src023[39] << 23) +
      (src023[40] << 23) +
      (src023[41] << 23) +
      (src023[42] << 23) +
      (src023[43] << 23) +
      (src023[44] << 23) +
      (src023[45] << 23) +
      (src023[46] << 23) +
      (src023[47] << 23) +
      (src023[48] << 23) +
      (src023[49] << 23) +
      (src023[50] << 23) +
      (src023[51] << 23) +
      (src023[52] << 23) +
      (src023[53] << 23) +
      (src023[54] << 23) +
      (src023[55] << 23) +
      (src023[56] << 23) +
      (src023[57] << 23) +
      (src023[58] << 23) +
      (src023[59] << 23) +
      (src023[60] << 23) +
      (src023[61] << 23) +
      (src023[62] << 23) +
      (src023[63] << 23) +
      (src023[64] << 23) +
      (src023[65] << 23) +
      (src023[66] << 23) +
      (src023[67] << 23) +
      (src023[68] << 23) +
      (src023[69] << 23) +
      (src023[70] << 23) +
      (src023[71] << 23) +
      (src023[72] << 23) +
      (src023[73] << 23) +
      (src023[74] << 23) +
      (src023[75] << 23) +
      (src023[76] << 23) +
      (src023[77] << 23) +
      (src023[78] << 23) +
      (src023[79] << 23) +
      (src023[80] << 23) +
      (src023[81] << 23) +
      (src023[82] << 23) +
      (src023[83] << 23) +
      (src023[84] << 23) +
      (src023[85] << 23) +
      (src023[86] << 23) +
      (src023[87] << 23) +
      (src023[88] << 23) +
      (src023[89] << 23) +
      (src023[90] << 23) +
      (src023[91] << 23) +
      (src023[92] << 23) +
      (src023[93] << 23) +
      (src023[94] << 23) +
      (src023[95] << 23) +
      (src023[96] << 23) +
      (src023[97] << 23) +
      (src023[98] << 23) +
      (src023[99] << 23) +
      (src023[100] << 23) +
      (src023[101] << 23) +
      (src023[102] << 23) +
      (src023[103] << 23) +
      (src023[104] << 23) +
      (src023[105] << 23) +
      (src023[106] << 23) +
      (src023[107] << 23) +
      (src023[108] << 23) +
      (src023[109] << 23) +
      (src023[110] << 23) +
      (src023[111] << 23) +
      (src023[112] << 23) +
      (src023[113] << 23) +
      (src023[114] << 23) +
      (src023[115] << 23) +
      (src023[116] << 23) +
      (src023[117] << 23) +
      (src023[118] << 23) +
      (src023[119] << 23) +
      (src023[120] << 23) +
      (src023[121] << 23) +
      (src023[122] << 23) +
      (src023[123] << 23) +
      (src023[124] << 23) +
      (src023[125] << 23) +
      (src023[126] << 23) +
      (src023[127] << 23) +
      (src024[0] << 24) +
      (src024[1] << 24) +
      (src024[2] << 24) +
      (src024[3] << 24) +
      (src024[4] << 24) +
      (src024[5] << 24) +
      (src024[6] << 24) +
      (src024[7] << 24) +
      (src024[8] << 24) +
      (src024[9] << 24) +
      (src024[10] << 24) +
      (src024[11] << 24) +
      (src024[12] << 24) +
      (src024[13] << 24) +
      (src024[14] << 24) +
      (src024[15] << 24) +
      (src024[16] << 24) +
      (src024[17] << 24) +
      (src024[18] << 24) +
      (src024[19] << 24) +
      (src024[20] << 24) +
      (src024[21] << 24) +
      (src024[22] << 24) +
      (src024[23] << 24) +
      (src024[24] << 24) +
      (src024[25] << 24) +
      (src024[26] << 24) +
      (src024[27] << 24) +
      (src024[28] << 24) +
      (src024[29] << 24) +
      (src024[30] << 24) +
      (src024[31] << 24) +
      (src024[32] << 24) +
      (src024[33] << 24) +
      (src024[34] << 24) +
      (src024[35] << 24) +
      (src024[36] << 24) +
      (src024[37] << 24) +
      (src024[38] << 24) +
      (src024[39] << 24) +
      (src024[40] << 24) +
      (src024[41] << 24) +
      (src024[42] << 24) +
      (src024[43] << 24) +
      (src024[44] << 24) +
      (src024[45] << 24) +
      (src024[46] << 24) +
      (src024[47] << 24) +
      (src024[48] << 24) +
      (src024[49] << 24) +
      (src024[50] << 24) +
      (src024[51] << 24) +
      (src024[52] << 24) +
      (src024[53] << 24) +
      (src024[54] << 24) +
      (src024[55] << 24) +
      (src024[56] << 24) +
      (src024[57] << 24) +
      (src024[58] << 24) +
      (src024[59] << 24) +
      (src024[60] << 24) +
      (src024[61] << 24) +
      (src024[62] << 24) +
      (src024[63] << 24) +
      (src024[64] << 24) +
      (src024[65] << 24) +
      (src024[66] << 24) +
      (src024[67] << 24) +
      (src024[68] << 24) +
      (src024[69] << 24) +
      (src024[70] << 24) +
      (src024[71] << 24) +
      (src024[72] << 24) +
      (src024[73] << 24) +
      (src024[74] << 24) +
      (src024[75] << 24) +
      (src024[76] << 24) +
      (src024[77] << 24) +
      (src024[78] << 24) +
      (src024[79] << 24) +
      (src024[80] << 24) +
      (src024[81] << 24) +
      (src024[82] << 24) +
      (src024[83] << 24) +
      (src024[84] << 24) +
      (src024[85] << 24) +
      (src024[86] << 24) +
      (src024[87] << 24) +
      (src024[88] << 24) +
      (src024[89] << 24) +
      (src024[90] << 24) +
      (src024[91] << 24) +
      (src024[92] << 24) +
      (src024[93] << 24) +
      (src024[94] << 24) +
      (src024[95] << 24) +
      (src024[96] << 24) +
      (src024[97] << 24) +
      (src024[98] << 24) +
      (src024[99] << 24) +
      (src024[100] << 24) +
      (src024[101] << 24) +
      (src024[102] << 24) +
      (src024[103] << 24) +
      (src024[104] << 24) +
      (src024[105] << 24) +
      (src024[106] << 24) +
      (src024[107] << 24) +
      (src024[108] << 24) +
      (src024[109] << 24) +
      (src024[110] << 24) +
      (src024[111] << 24) +
      (src024[112] << 24) +
      (src024[113] << 24) +
      (src024[114] << 24) +
      (src024[115] << 24) +
      (src024[116] << 24) +
      (src024[117] << 24) +
      (src024[118] << 24) +
      (src024[119] << 24) +
      (src024[120] << 24) +
      (src024[121] << 24) +
      (src024[122] << 24) +
      (src024[123] << 24) +
      (src024[124] << 24) +
      (src024[125] << 24) +
      (src024[126] << 24) +
      (src024[127] << 24) +
      (src025[0] << 25) +
      (src025[1] << 25) +
      (src025[2] << 25) +
      (src025[3] << 25) +
      (src025[4] << 25) +
      (src025[5] << 25) +
      (src025[6] << 25) +
      (src025[7] << 25) +
      (src025[8] << 25) +
      (src025[9] << 25) +
      (src025[10] << 25) +
      (src025[11] << 25) +
      (src025[12] << 25) +
      (src025[13] << 25) +
      (src025[14] << 25) +
      (src025[15] << 25) +
      (src025[16] << 25) +
      (src025[17] << 25) +
      (src025[18] << 25) +
      (src025[19] << 25) +
      (src025[20] << 25) +
      (src025[21] << 25) +
      (src025[22] << 25) +
      (src025[23] << 25) +
      (src025[24] << 25) +
      (src025[25] << 25) +
      (src025[26] << 25) +
      (src025[27] << 25) +
      (src025[28] << 25) +
      (src025[29] << 25) +
      (src025[30] << 25) +
      (src025[31] << 25) +
      (src025[32] << 25) +
      (src025[33] << 25) +
      (src025[34] << 25) +
      (src025[35] << 25) +
      (src025[36] << 25) +
      (src025[37] << 25) +
      (src025[38] << 25) +
      (src025[39] << 25) +
      (src025[40] << 25) +
      (src025[41] << 25) +
      (src025[42] << 25) +
      (src025[43] << 25) +
      (src025[44] << 25) +
      (src025[45] << 25) +
      (src025[46] << 25) +
      (src025[47] << 25) +
      (src025[48] << 25) +
      (src025[49] << 25) +
      (src025[50] << 25) +
      (src025[51] << 25) +
      (src025[52] << 25) +
      (src025[53] << 25) +
      (src025[54] << 25) +
      (src025[55] << 25) +
      (src025[56] << 25) +
      (src025[57] << 25) +
      (src025[58] << 25) +
      (src025[59] << 25) +
      (src025[60] << 25) +
      (src025[61] << 25) +
      (src025[62] << 25) +
      (src025[63] << 25) +
      (src025[64] << 25) +
      (src025[65] << 25) +
      (src025[66] << 25) +
      (src025[67] << 25) +
      (src025[68] << 25) +
      (src025[69] << 25) +
      (src025[70] << 25) +
      (src025[71] << 25) +
      (src025[72] << 25) +
      (src025[73] << 25) +
      (src025[74] << 25) +
      (src025[75] << 25) +
      (src025[76] << 25) +
      (src025[77] << 25) +
      (src025[78] << 25) +
      (src025[79] << 25) +
      (src025[80] << 25) +
      (src025[81] << 25) +
      (src025[82] << 25) +
      (src025[83] << 25) +
      (src025[84] << 25) +
      (src025[85] << 25) +
      (src025[86] << 25) +
      (src025[87] << 25) +
      (src025[88] << 25) +
      (src025[89] << 25) +
      (src025[90] << 25) +
      (src025[91] << 25) +
      (src025[92] << 25) +
      (src025[93] << 25) +
      (src025[94] << 25) +
      (src025[95] << 25) +
      (src025[96] << 25) +
      (src025[97] << 25) +
      (src025[98] << 25) +
      (src025[99] << 25) +
      (src025[100] << 25) +
      (src025[101] << 25) +
      (src025[102] << 25) +
      (src025[103] << 25) +
      (src025[104] << 25) +
      (src025[105] << 25) +
      (src025[106] << 25) +
      (src025[107] << 25) +
      (src025[108] << 25) +
      (src025[109] << 25) +
      (src025[110] << 25) +
      (src025[111] << 25) +
      (src025[112] << 25) +
      (src025[113] << 25) +
      (src025[114] << 25) +
      (src025[115] << 25) +
      (src025[116] << 25) +
      (src025[117] << 25) +
      (src025[118] << 25) +
      (src025[119] << 25) +
      (src025[120] << 25) +
      (src025[121] << 25) +
      (src025[122] << 25) +
      (src025[123] << 25) +
      (src025[124] << 25) +
      (src025[125] << 25) +
      (src025[126] << 25) +
      (src025[127] << 25) +
      (src026[0] << 26) +
      (src026[1] << 26) +
      (src026[2] << 26) +
      (src026[3] << 26) +
      (src026[4] << 26) +
      (src026[5] << 26) +
      (src026[6] << 26) +
      (src026[7] << 26) +
      (src026[8] << 26) +
      (src026[9] << 26) +
      (src026[10] << 26) +
      (src026[11] << 26) +
      (src026[12] << 26) +
      (src026[13] << 26) +
      (src026[14] << 26) +
      (src026[15] << 26) +
      (src026[16] << 26) +
      (src026[17] << 26) +
      (src026[18] << 26) +
      (src026[19] << 26) +
      (src026[20] << 26) +
      (src026[21] << 26) +
      (src026[22] << 26) +
      (src026[23] << 26) +
      (src026[24] << 26) +
      (src026[25] << 26) +
      (src026[26] << 26) +
      (src026[27] << 26) +
      (src026[28] << 26) +
      (src026[29] << 26) +
      (src026[30] << 26) +
      (src026[31] << 26) +
      (src026[32] << 26) +
      (src026[33] << 26) +
      (src026[34] << 26) +
      (src026[35] << 26) +
      (src026[36] << 26) +
      (src026[37] << 26) +
      (src026[38] << 26) +
      (src026[39] << 26) +
      (src026[40] << 26) +
      (src026[41] << 26) +
      (src026[42] << 26) +
      (src026[43] << 26) +
      (src026[44] << 26) +
      (src026[45] << 26) +
      (src026[46] << 26) +
      (src026[47] << 26) +
      (src026[48] << 26) +
      (src026[49] << 26) +
      (src026[50] << 26) +
      (src026[51] << 26) +
      (src026[52] << 26) +
      (src026[53] << 26) +
      (src026[54] << 26) +
      (src026[55] << 26) +
      (src026[56] << 26) +
      (src026[57] << 26) +
      (src026[58] << 26) +
      (src026[59] << 26) +
      (src026[60] << 26) +
      (src026[61] << 26) +
      (src026[62] << 26) +
      (src026[63] << 26) +
      (src026[64] << 26) +
      (src026[65] << 26) +
      (src026[66] << 26) +
      (src026[67] << 26) +
      (src026[68] << 26) +
      (src026[69] << 26) +
      (src026[70] << 26) +
      (src026[71] << 26) +
      (src026[72] << 26) +
      (src026[73] << 26) +
      (src026[74] << 26) +
      (src026[75] << 26) +
      (src026[76] << 26) +
      (src026[77] << 26) +
      (src026[78] << 26) +
      (src026[79] << 26) +
      (src026[80] << 26) +
      (src026[81] << 26) +
      (src026[82] << 26) +
      (src026[83] << 26) +
      (src026[84] << 26) +
      (src026[85] << 26) +
      (src026[86] << 26) +
      (src026[87] << 26) +
      (src026[88] << 26) +
      (src026[89] << 26) +
      (src026[90] << 26) +
      (src026[91] << 26) +
      (src026[92] << 26) +
      (src026[93] << 26) +
      (src026[94] << 26) +
      (src026[95] << 26) +
      (src026[96] << 26) +
      (src026[97] << 26) +
      (src026[98] << 26) +
      (src026[99] << 26) +
      (src026[100] << 26) +
      (src026[101] << 26) +
      (src026[102] << 26) +
      (src026[103] << 26) +
      (src026[104] << 26) +
      (src026[105] << 26) +
      (src026[106] << 26) +
      (src026[107] << 26) +
      (src026[108] << 26) +
      (src026[109] << 26) +
      (src026[110] << 26) +
      (src026[111] << 26) +
      (src026[112] << 26) +
      (src026[113] << 26) +
      (src026[114] << 26) +
      (src026[115] << 26) +
      (src026[116] << 26) +
      (src026[117] << 26) +
      (src026[118] << 26) +
      (src026[119] << 26) +
      (src026[120] << 26) +
      (src026[121] << 26) +
      (src026[122] << 26) +
      (src026[123] << 26) +
      (src026[124] << 26) +
      (src026[125] << 26) +
      (src026[126] << 26) +
      (src026[127] << 26) +
      (src027[0] << 27) +
      (src027[1] << 27) +
      (src027[2] << 27) +
      (src027[3] << 27) +
      (src027[4] << 27) +
      (src027[5] << 27) +
      (src027[6] << 27) +
      (src027[7] << 27) +
      (src027[8] << 27) +
      (src027[9] << 27) +
      (src027[10] << 27) +
      (src027[11] << 27) +
      (src027[12] << 27) +
      (src027[13] << 27) +
      (src027[14] << 27) +
      (src027[15] << 27) +
      (src027[16] << 27) +
      (src027[17] << 27) +
      (src027[18] << 27) +
      (src027[19] << 27) +
      (src027[20] << 27) +
      (src027[21] << 27) +
      (src027[22] << 27) +
      (src027[23] << 27) +
      (src027[24] << 27) +
      (src027[25] << 27) +
      (src027[26] << 27) +
      (src027[27] << 27) +
      (src027[28] << 27) +
      (src027[29] << 27) +
      (src027[30] << 27) +
      (src027[31] << 27) +
      (src027[32] << 27) +
      (src027[33] << 27) +
      (src027[34] << 27) +
      (src027[35] << 27) +
      (src027[36] << 27) +
      (src027[37] << 27) +
      (src027[38] << 27) +
      (src027[39] << 27) +
      (src027[40] << 27) +
      (src027[41] << 27) +
      (src027[42] << 27) +
      (src027[43] << 27) +
      (src027[44] << 27) +
      (src027[45] << 27) +
      (src027[46] << 27) +
      (src027[47] << 27) +
      (src027[48] << 27) +
      (src027[49] << 27) +
      (src027[50] << 27) +
      (src027[51] << 27) +
      (src027[52] << 27) +
      (src027[53] << 27) +
      (src027[54] << 27) +
      (src027[55] << 27) +
      (src027[56] << 27) +
      (src027[57] << 27) +
      (src027[58] << 27) +
      (src027[59] << 27) +
      (src027[60] << 27) +
      (src027[61] << 27) +
      (src027[62] << 27) +
      (src027[63] << 27) +
      (src027[64] << 27) +
      (src027[65] << 27) +
      (src027[66] << 27) +
      (src027[67] << 27) +
      (src027[68] << 27) +
      (src027[69] << 27) +
      (src027[70] << 27) +
      (src027[71] << 27) +
      (src027[72] << 27) +
      (src027[73] << 27) +
      (src027[74] << 27) +
      (src027[75] << 27) +
      (src027[76] << 27) +
      (src027[77] << 27) +
      (src027[78] << 27) +
      (src027[79] << 27) +
      (src027[80] << 27) +
      (src027[81] << 27) +
      (src027[82] << 27) +
      (src027[83] << 27) +
      (src027[84] << 27) +
      (src027[85] << 27) +
      (src027[86] << 27) +
      (src027[87] << 27) +
      (src027[88] << 27) +
      (src027[89] << 27) +
      (src027[90] << 27) +
      (src027[91] << 27) +
      (src027[92] << 27) +
      (src027[93] << 27) +
      (src027[94] << 27) +
      (src027[95] << 27) +
      (src027[96] << 27) +
      (src027[97] << 27) +
      (src027[98] << 27) +
      (src027[99] << 27) +
      (src027[100] << 27) +
      (src027[101] << 27) +
      (src027[102] << 27) +
      (src027[103] << 27) +
      (src027[104] << 27) +
      (src027[105] << 27) +
      (src027[106] << 27) +
      (src027[107] << 27) +
      (src027[108] << 27) +
      (src027[109] << 27) +
      (src027[110] << 27) +
      (src027[111] << 27) +
      (src027[112] << 27) +
      (src027[113] << 27) +
      (src027[114] << 27) +
      (src027[115] << 27) +
      (src027[116] << 27) +
      (src027[117] << 27) +
      (src027[118] << 27) +
      (src027[119] << 27) +
      (src027[120] << 27) +
      (src027[121] << 27) +
      (src027[122] << 27) +
      (src027[123] << 27) +
      (src027[124] << 27) +
      (src027[125] << 27) +
      (src027[126] << 27) +
      (src027[127] << 27) +
      (src028[0] << 28) +
      (src028[1] << 28) +
      (src028[2] << 28) +
      (src028[3] << 28) +
      (src028[4] << 28) +
      (src028[5] << 28) +
      (src028[6] << 28) +
      (src028[7] << 28) +
      (src028[8] << 28) +
      (src028[9] << 28) +
      (src028[10] << 28) +
      (src028[11] << 28) +
      (src028[12] << 28) +
      (src028[13] << 28) +
      (src028[14] << 28) +
      (src028[15] << 28) +
      (src028[16] << 28) +
      (src028[17] << 28) +
      (src028[18] << 28) +
      (src028[19] << 28) +
      (src028[20] << 28) +
      (src028[21] << 28) +
      (src028[22] << 28) +
      (src028[23] << 28) +
      (src028[24] << 28) +
      (src028[25] << 28) +
      (src028[26] << 28) +
      (src028[27] << 28) +
      (src028[28] << 28) +
      (src028[29] << 28) +
      (src028[30] << 28) +
      (src028[31] << 28) +
      (src028[32] << 28) +
      (src028[33] << 28) +
      (src028[34] << 28) +
      (src028[35] << 28) +
      (src028[36] << 28) +
      (src028[37] << 28) +
      (src028[38] << 28) +
      (src028[39] << 28) +
      (src028[40] << 28) +
      (src028[41] << 28) +
      (src028[42] << 28) +
      (src028[43] << 28) +
      (src028[44] << 28) +
      (src028[45] << 28) +
      (src028[46] << 28) +
      (src028[47] << 28) +
      (src028[48] << 28) +
      (src028[49] << 28) +
      (src028[50] << 28) +
      (src028[51] << 28) +
      (src028[52] << 28) +
      (src028[53] << 28) +
      (src028[54] << 28) +
      (src028[55] << 28) +
      (src028[56] << 28) +
      (src028[57] << 28) +
      (src028[58] << 28) +
      (src028[59] << 28) +
      (src028[60] << 28) +
      (src028[61] << 28) +
      (src028[62] << 28) +
      (src028[63] << 28) +
      (src028[64] << 28) +
      (src028[65] << 28) +
      (src028[66] << 28) +
      (src028[67] << 28) +
      (src028[68] << 28) +
      (src028[69] << 28) +
      (src028[70] << 28) +
      (src028[71] << 28) +
      (src028[72] << 28) +
      (src028[73] << 28) +
      (src028[74] << 28) +
      (src028[75] << 28) +
      (src028[76] << 28) +
      (src028[77] << 28) +
      (src028[78] << 28) +
      (src028[79] << 28) +
      (src028[80] << 28) +
      (src028[81] << 28) +
      (src028[82] << 28) +
      (src028[83] << 28) +
      (src028[84] << 28) +
      (src028[85] << 28) +
      (src028[86] << 28) +
      (src028[87] << 28) +
      (src028[88] << 28) +
      (src028[89] << 28) +
      (src028[90] << 28) +
      (src028[91] << 28) +
      (src028[92] << 28) +
      (src028[93] << 28) +
      (src028[94] << 28) +
      (src028[95] << 28) +
      (src028[96] << 28) +
      (src028[97] << 28) +
      (src028[98] << 28) +
      (src028[99] << 28) +
      (src028[100] << 28) +
      (src028[101] << 28) +
      (src028[102] << 28) +
      (src028[103] << 28) +
      (src028[104] << 28) +
      (src028[105] << 28) +
      (src028[106] << 28) +
      (src028[107] << 28) +
      (src028[108] << 28) +
      (src028[109] << 28) +
      (src028[110] << 28) +
      (src028[111] << 28) +
      (src028[112] << 28) +
      (src028[113] << 28) +
      (src028[114] << 28) +
      (src028[115] << 28) +
      (src028[116] << 28) +
      (src028[117] << 28) +
      (src028[118] << 28) +
      (src028[119] << 28) +
      (src028[120] << 28) +
      (src028[121] << 28) +
      (src028[122] << 28) +
      (src028[123] << 28) +
      (src028[124] << 28) +
      (src028[125] << 28) +
      (src028[126] << 28) +
      (src028[127] << 28) +
      (src029[0] << 29) +
      (src029[1] << 29) +
      (src029[2] << 29) +
      (src029[3] << 29) +
      (src029[4] << 29) +
      (src029[5] << 29) +
      (src029[6] << 29) +
      (src029[7] << 29) +
      (src029[8] << 29) +
      (src029[9] << 29) +
      (src029[10] << 29) +
      (src029[11] << 29) +
      (src029[12] << 29) +
      (src029[13] << 29) +
      (src029[14] << 29) +
      (src029[15] << 29) +
      (src029[16] << 29) +
      (src029[17] << 29) +
      (src029[18] << 29) +
      (src029[19] << 29) +
      (src029[20] << 29) +
      (src029[21] << 29) +
      (src029[22] << 29) +
      (src029[23] << 29) +
      (src029[24] << 29) +
      (src029[25] << 29) +
      (src029[26] << 29) +
      (src029[27] << 29) +
      (src029[28] << 29) +
      (src029[29] << 29) +
      (src029[30] << 29) +
      (src029[31] << 29) +
      (src029[32] << 29) +
      (src029[33] << 29) +
      (src029[34] << 29) +
      (src029[35] << 29) +
      (src029[36] << 29) +
      (src029[37] << 29) +
      (src029[38] << 29) +
      (src029[39] << 29) +
      (src029[40] << 29) +
      (src029[41] << 29) +
      (src029[42] << 29) +
      (src029[43] << 29) +
      (src029[44] << 29) +
      (src029[45] << 29) +
      (src029[46] << 29) +
      (src029[47] << 29) +
      (src029[48] << 29) +
      (src029[49] << 29) +
      (src029[50] << 29) +
      (src029[51] << 29) +
      (src029[52] << 29) +
      (src029[53] << 29) +
      (src029[54] << 29) +
      (src029[55] << 29) +
      (src029[56] << 29) +
      (src029[57] << 29) +
      (src029[58] << 29) +
      (src029[59] << 29) +
      (src029[60] << 29) +
      (src029[61] << 29) +
      (src029[62] << 29) +
      (src029[63] << 29) +
      (src029[64] << 29) +
      (src029[65] << 29) +
      (src029[66] << 29) +
      (src029[67] << 29) +
      (src029[68] << 29) +
      (src029[69] << 29) +
      (src029[70] << 29) +
      (src029[71] << 29) +
      (src029[72] << 29) +
      (src029[73] << 29) +
      (src029[74] << 29) +
      (src029[75] << 29) +
      (src029[76] << 29) +
      (src029[77] << 29) +
      (src029[78] << 29) +
      (src029[79] << 29) +
      (src029[80] << 29) +
      (src029[81] << 29) +
      (src029[82] << 29) +
      (src029[83] << 29) +
      (src029[84] << 29) +
      (src029[85] << 29) +
      (src029[86] << 29) +
      (src029[87] << 29) +
      (src029[88] << 29) +
      (src029[89] << 29) +
      (src029[90] << 29) +
      (src029[91] << 29) +
      (src029[92] << 29) +
      (src029[93] << 29) +
      (src029[94] << 29) +
      (src029[95] << 29) +
      (src029[96] << 29) +
      (src029[97] << 29) +
      (src029[98] << 29) +
      (src029[99] << 29) +
      (src029[100] << 29) +
      (src029[101] << 29) +
      (src029[102] << 29) +
      (src029[103] << 29) +
      (src029[104] << 29) +
      (src029[105] << 29) +
      (src029[106] << 29) +
      (src029[107] << 29) +
      (src029[108] << 29) +
      (src029[109] << 29) +
      (src029[110] << 29) +
      (src029[111] << 29) +
      (src029[112] << 29) +
      (src029[113] << 29) +
      (src029[114] << 29) +
      (src029[115] << 29) +
      (src029[116] << 29) +
      (src029[117] << 29) +
      (src029[118] << 29) +
      (src029[119] << 29) +
      (src029[120] << 29) +
      (src029[121] << 29) +
      (src029[122] << 29) +
      (src029[123] << 29) +
      (src029[124] << 29) +
      (src029[125] << 29) +
      (src029[126] << 29) +
      (src029[127] << 29) +
      (src030[0] << 30) +
      (src030[1] << 30) +
      (src030[2] << 30) +
      (src030[3] << 30) +
      (src030[4] << 30) +
      (src030[5] << 30) +
      (src030[6] << 30) +
      (src030[7] << 30) +
      (src030[8] << 30) +
      (src030[9] << 30) +
      (src030[10] << 30) +
      (src030[11] << 30) +
      (src030[12] << 30) +
      (src030[13] << 30) +
      (src030[14] << 30) +
      (src030[15] << 30) +
      (src030[16] << 30) +
      (src030[17] << 30) +
      (src030[18] << 30) +
      (src030[19] << 30) +
      (src030[20] << 30) +
      (src030[21] << 30) +
      (src030[22] << 30) +
      (src030[23] << 30) +
      (src030[24] << 30) +
      (src030[25] << 30) +
      (src030[26] << 30) +
      (src030[27] << 30) +
      (src030[28] << 30) +
      (src030[29] << 30) +
      (src030[30] << 30) +
      (src030[31] << 30) +
      (src030[32] << 30) +
      (src030[33] << 30) +
      (src030[34] << 30) +
      (src030[35] << 30) +
      (src030[36] << 30) +
      (src030[37] << 30) +
      (src030[38] << 30) +
      (src030[39] << 30) +
      (src030[40] << 30) +
      (src030[41] << 30) +
      (src030[42] << 30) +
      (src030[43] << 30) +
      (src030[44] << 30) +
      (src030[45] << 30) +
      (src030[46] << 30) +
      (src030[47] << 30) +
      (src030[48] << 30) +
      (src030[49] << 30) +
      (src030[50] << 30) +
      (src030[51] << 30) +
      (src030[52] << 30) +
      (src030[53] << 30) +
      (src030[54] << 30) +
      (src030[55] << 30) +
      (src030[56] << 30) +
      (src030[57] << 30) +
      (src030[58] << 30) +
      (src030[59] << 30) +
      (src030[60] << 30) +
      (src030[61] << 30) +
      (src030[62] << 30) +
      (src030[63] << 30) +
      (src030[64] << 30) +
      (src030[65] << 30) +
      (src030[66] << 30) +
      (src030[67] << 30) +
      (src030[68] << 30) +
      (src030[69] << 30) +
      (src030[70] << 30) +
      (src030[71] << 30) +
      (src030[72] << 30) +
      (src030[73] << 30) +
      (src030[74] << 30) +
      (src030[75] << 30) +
      (src030[76] << 30) +
      (src030[77] << 30) +
      (src030[78] << 30) +
      (src030[79] << 30) +
      (src030[80] << 30) +
      (src030[81] << 30) +
      (src030[82] << 30) +
      (src030[83] << 30) +
      (src030[84] << 30) +
      (src030[85] << 30) +
      (src030[86] << 30) +
      (src030[87] << 30) +
      (src030[88] << 30) +
      (src030[89] << 30) +
      (src030[90] << 30) +
      (src030[91] << 30) +
      (src030[92] << 30) +
      (src030[93] << 30) +
      (src030[94] << 30) +
      (src030[95] << 30) +
      (src030[96] << 30) +
      (src030[97] << 30) +
      (src030[98] << 30) +
      (src030[99] << 30) +
      (src030[100] << 30) +
      (src030[101] << 30) +
      (src030[102] << 30) +
      (src030[103] << 30) +
      (src030[104] << 30) +
      (src030[105] << 30) +
      (src030[106] << 30) +
      (src030[107] << 30) +
      (src030[108] << 30) +
      (src030[109] << 30) +
      (src030[110] << 30) +
      (src030[111] << 30) +
      (src030[112] << 30) +
      (src030[113] << 30) +
      (src030[114] << 30) +
      (src030[115] << 30) +
      (src030[116] << 30) +
      (src030[117] << 30) +
      (src030[118] << 30) +
      (src030[119] << 30) +
      (src030[120] << 30) +
      (src030[121] << 30) +
      (src030[122] << 30) +
      (src030[123] << 30) +
      (src030[124] << 30) +
      (src030[125] << 30) +
      (src030[126] << 30) +
      (src030[127] << 30) +
      (src031[0] << 31) +
      (src031[1] << 31) +
      (src031[2] << 31) +
      (src031[3] << 31) +
      (src031[4] << 31) +
      (src031[5] << 31) +
      (src031[6] << 31) +
      (src031[7] << 31) +
      (src031[8] << 31) +
      (src031[9] << 31) +
      (src031[10] << 31) +
      (src031[11] << 31) +
      (src031[12] << 31) +
      (src031[13] << 31) +
      (src031[14] << 31) +
      (src031[15] << 31) +
      (src031[16] << 31) +
      (src031[17] << 31) +
      (src031[18] << 31) +
      (src031[19] << 31) +
      (src031[20] << 31) +
      (src031[21] << 31) +
      (src031[22] << 31) +
      (src031[23] << 31) +
      (src031[24] << 31) +
      (src031[25] << 31) +
      (src031[26] << 31) +
      (src031[27] << 31) +
      (src031[28] << 31) +
      (src031[29] << 31) +
      (src031[30] << 31) +
      (src031[31] << 31) +
      (src031[32] << 31) +
      (src031[33] << 31) +
      (src031[34] << 31) +
      (src031[35] << 31) +
      (src031[36] << 31) +
      (src031[37] << 31) +
      (src031[38] << 31) +
      (src031[39] << 31) +
      (src031[40] << 31) +
      (src031[41] << 31) +
      (src031[42] << 31) +
      (src031[43] << 31) +
      (src031[44] << 31) +
      (src031[45] << 31) +
      (src031[46] << 31) +
      (src031[47] << 31) +
      (src031[48] << 31) +
      (src031[49] << 31) +
      (src031[50] << 31) +
      (src031[51] << 31) +
      (src031[52] << 31) +
      (src031[53] << 31) +
      (src031[54] << 31) +
      (src031[55] << 31) +
      (src031[56] << 31) +
      (src031[57] << 31) +
      (src031[58] << 31) +
      (src031[59] << 31) +
      (src031[60] << 31) +
      (src031[61] << 31) +
      (src031[62] << 31) +
      (src031[63] << 31) +
      (src031[64] << 31) +
      (src031[65] << 31) +
      (src031[66] << 31) +
      (src031[67] << 31) +
      (src031[68] << 31) +
      (src031[69] << 31) +
      (src031[70] << 31) +
      (src031[71] << 31) +
      (src031[72] << 31) +
      (src031[73] << 31) +
      (src031[74] << 31) +
      (src031[75] << 31) +
      (src031[76] << 31) +
      (src031[77] << 31) +
      (src031[78] << 31) +
      (src031[79] << 31) +
      (src031[80] << 31) +
      (src031[81] << 31) +
      (src031[82] << 31) +
      (src031[83] << 31) +
      (src031[84] << 31) +
      (src031[85] << 31) +
      (src031[86] << 31) +
      (src031[87] << 31) +
      (src031[88] << 31) +
      (src031[89] << 31) +
      (src031[90] << 31) +
      (src031[91] << 31) +
      (src031[92] << 31) +
      (src031[93] << 31) +
      (src031[94] << 31) +
      (src031[95] << 31) +
      (src031[96] << 31) +
      (src031[97] << 31) +
      (src031[98] << 31) +
      (src031[99] << 31) +
      (src031[100] << 31) +
      (src031[101] << 31) +
      (src031[102] << 31) +
      (src031[103] << 31) +
      (src031[104] << 31) +
      (src031[105] << 31) +
      (src031[106] << 31) +
      (src031[107] << 31) +
      (src031[108] << 31) +
      (src031[109] << 31) +
      (src031[110] << 31) +
      (src031[111] << 31) +
      (src031[112] << 31) +
      (src031[113] << 31) +
      (src031[114] << 31) +
      (src031[115] << 31) +
      (src031[116] << 31) +
      (src031[117] << 31) +
      (src031[118] << 31) +
      (src031[119] << 31) +
      (src031[120] << 31) +
      (src031[121] << 31) +
      (src031[122] << 31) +
      (src031[123] << 31) +
      (src031[124] << 31) +
      (src031[125] << 31) +
      (src031[126] << 31) +
      (src031[127] << 31) +
      (src032[0] << 32) +
      (src032[1] << 32) +
      (src032[2] << 32) +
      (src032[3] << 32) +
      (src032[4] << 32) +
      (src032[5] << 32) +
      (src032[6] << 32) +
      (src032[7] << 32) +
      (src032[8] << 32) +
      (src032[9] << 32) +
      (src032[10] << 32) +
      (src032[11] << 32) +
      (src032[12] << 32) +
      (src032[13] << 32) +
      (src032[14] << 32) +
      (src032[15] << 32) +
      (src032[16] << 32) +
      (src032[17] << 32) +
      (src032[18] << 32) +
      (src032[19] << 32) +
      (src032[20] << 32) +
      (src032[21] << 32) +
      (src032[22] << 32) +
      (src032[23] << 32) +
      (src032[24] << 32) +
      (src032[25] << 32) +
      (src032[26] << 32) +
      (src032[27] << 32) +
      (src032[28] << 32) +
      (src032[29] << 32) +
      (src032[30] << 32) +
      (src032[31] << 32) +
      (src032[32] << 32) +
      (src032[33] << 32) +
      (src032[34] << 32) +
      (src032[35] << 32) +
      (src032[36] << 32) +
      (src032[37] << 32) +
      (src032[38] << 32) +
      (src032[39] << 32) +
      (src032[40] << 32) +
      (src032[41] << 32) +
      (src032[42] << 32) +
      (src032[43] << 32) +
      (src032[44] << 32) +
      (src032[45] << 32) +
      (src032[46] << 32) +
      (src032[47] << 32) +
      (src032[48] << 32) +
      (src032[49] << 32) +
      (src032[50] << 32) +
      (src032[51] << 32) +
      (src032[52] << 32) +
      (src032[53] << 32) +
      (src032[54] << 32) +
      (src032[55] << 32) +
      (src032[56] << 32) +
      (src032[57] << 32) +
      (src032[58] << 32) +
      (src032[59] << 32) +
      (src032[60] << 32) +
      (src032[61] << 32) +
      (src032[62] << 32) +
      (src032[63] << 32) +
      (src032[64] << 32) +
      (src032[65] << 32) +
      (src032[66] << 32) +
      (src032[67] << 32) +
      (src032[68] << 32) +
      (src032[69] << 32) +
      (src032[70] << 32) +
      (src032[71] << 32) +
      (src032[72] << 32) +
      (src032[73] << 32) +
      (src032[74] << 32) +
      (src032[75] << 32) +
      (src032[76] << 32) +
      (src032[77] << 32) +
      (src032[78] << 32) +
      (src032[79] << 32) +
      (src032[80] << 32) +
      (src032[81] << 32) +
      (src032[82] << 32) +
      (src032[83] << 32) +
      (src032[84] << 32) +
      (src032[85] << 32) +
      (src032[86] << 32) +
      (src032[87] << 32) +
      (src032[88] << 32) +
      (src032[89] << 32) +
      (src032[90] << 32) +
      (src032[91] << 32) +
      (src032[92] << 32) +
      (src032[93] << 32) +
      (src032[94] << 32) +
      (src032[95] << 32) +
      (src032[96] << 32) +
      (src032[97] << 32) +
      (src032[98] << 32) +
      (src032[99] << 32) +
      (src032[100] << 32) +
      (src032[101] << 32) +
      (src032[102] << 32) +
      (src032[103] << 32) +
      (src032[104] << 32) +
      (src032[105] << 32) +
      (src032[106] << 32) +
      (src032[107] << 32) +
      (src032[108] << 32) +
      (src032[109] << 32) +
      (src032[110] << 32) +
      (src032[111] << 32) +
      (src032[112] << 32) +
      (src032[113] << 32) +
      (src032[114] << 32) +
      (src032[115] << 32) +
      (src032[116] << 32) +
      (src032[117] << 32) +
      (src032[118] << 32) +
      (src032[119] << 32) +
      (src032[120] << 32) +
      (src032[121] << 32) +
      (src032[122] << 32) +
      (src032[123] << 32) +
      (src032[124] << 32) +
      (src032[125] << 32) +
      (src032[126] << 32) +
      (src032[127] << 32) +
      (src033[0] << 33) +
      (src033[1] << 33) +
      (src033[2] << 33) +
      (src033[3] << 33) +
      (src033[4] << 33) +
      (src033[5] << 33) +
      (src033[6] << 33) +
      (src033[7] << 33) +
      (src033[8] << 33) +
      (src033[9] << 33) +
      (src033[10] << 33) +
      (src033[11] << 33) +
      (src033[12] << 33) +
      (src033[13] << 33) +
      (src033[14] << 33) +
      (src033[15] << 33) +
      (src033[16] << 33) +
      (src033[17] << 33) +
      (src033[18] << 33) +
      (src033[19] << 33) +
      (src033[20] << 33) +
      (src033[21] << 33) +
      (src033[22] << 33) +
      (src033[23] << 33) +
      (src033[24] << 33) +
      (src033[25] << 33) +
      (src033[26] << 33) +
      (src033[27] << 33) +
      (src033[28] << 33) +
      (src033[29] << 33) +
      (src033[30] << 33) +
      (src033[31] << 33) +
      (src033[32] << 33) +
      (src033[33] << 33) +
      (src033[34] << 33) +
      (src033[35] << 33) +
      (src033[36] << 33) +
      (src033[37] << 33) +
      (src033[38] << 33) +
      (src033[39] << 33) +
      (src033[40] << 33) +
      (src033[41] << 33) +
      (src033[42] << 33) +
      (src033[43] << 33) +
      (src033[44] << 33) +
      (src033[45] << 33) +
      (src033[46] << 33) +
      (src033[47] << 33) +
      (src033[48] << 33) +
      (src033[49] << 33) +
      (src033[50] << 33) +
      (src033[51] << 33) +
      (src033[52] << 33) +
      (src033[53] << 33) +
      (src033[54] << 33) +
      (src033[55] << 33) +
      (src033[56] << 33) +
      (src033[57] << 33) +
      (src033[58] << 33) +
      (src033[59] << 33) +
      (src033[60] << 33) +
      (src033[61] << 33) +
      (src033[62] << 33) +
      (src033[63] << 33) +
      (src033[64] << 33) +
      (src033[65] << 33) +
      (src033[66] << 33) +
      (src033[67] << 33) +
      (src033[68] << 33) +
      (src033[69] << 33) +
      (src033[70] << 33) +
      (src033[71] << 33) +
      (src033[72] << 33) +
      (src033[73] << 33) +
      (src033[74] << 33) +
      (src033[75] << 33) +
      (src033[76] << 33) +
      (src033[77] << 33) +
      (src033[78] << 33) +
      (src033[79] << 33) +
      (src033[80] << 33) +
      (src033[81] << 33) +
      (src033[82] << 33) +
      (src033[83] << 33) +
      (src033[84] << 33) +
      (src033[85] << 33) +
      (src033[86] << 33) +
      (src033[87] << 33) +
      (src033[88] << 33) +
      (src033[89] << 33) +
      (src033[90] << 33) +
      (src033[91] << 33) +
      (src033[92] << 33) +
      (src033[93] << 33) +
      (src033[94] << 33) +
      (src033[95] << 33) +
      (src033[96] << 33) +
      (src033[97] << 33) +
      (src033[98] << 33) +
      (src033[99] << 33) +
      (src033[100] << 33) +
      (src033[101] << 33) +
      (src033[102] << 33) +
      (src033[103] << 33) +
      (src033[104] << 33) +
      (src033[105] << 33) +
      (src033[106] << 33) +
      (src033[107] << 33) +
      (src033[108] << 33) +
      (src033[109] << 33) +
      (src033[110] << 33) +
      (src033[111] << 33) +
      (src033[112] << 33) +
      (src033[113] << 33) +
      (src033[114] << 33) +
      (src033[115] << 33) +
      (src033[116] << 33) +
      (src033[117] << 33) +
      (src033[118] << 33) +
      (src033[119] << 33) +
      (src033[120] << 33) +
      (src033[121] << 33) +
      (src033[122] << 33) +
      (src033[123] << 33) +
      (src033[124] << 33) +
      (src033[125] << 33) +
      (src033[126] << 33) +
      (src033[127] << 33) +
      (src034[0] << 34) +
      (src034[1] << 34) +
      (src034[2] << 34) +
      (src034[3] << 34) +
      (src034[4] << 34) +
      (src034[5] << 34) +
      (src034[6] << 34) +
      (src034[7] << 34) +
      (src034[8] << 34) +
      (src034[9] << 34) +
      (src034[10] << 34) +
      (src034[11] << 34) +
      (src034[12] << 34) +
      (src034[13] << 34) +
      (src034[14] << 34) +
      (src034[15] << 34) +
      (src034[16] << 34) +
      (src034[17] << 34) +
      (src034[18] << 34) +
      (src034[19] << 34) +
      (src034[20] << 34) +
      (src034[21] << 34) +
      (src034[22] << 34) +
      (src034[23] << 34) +
      (src034[24] << 34) +
      (src034[25] << 34) +
      (src034[26] << 34) +
      (src034[27] << 34) +
      (src034[28] << 34) +
      (src034[29] << 34) +
      (src034[30] << 34) +
      (src034[31] << 34) +
      (src034[32] << 34) +
      (src034[33] << 34) +
      (src034[34] << 34) +
      (src034[35] << 34) +
      (src034[36] << 34) +
      (src034[37] << 34) +
      (src034[38] << 34) +
      (src034[39] << 34) +
      (src034[40] << 34) +
      (src034[41] << 34) +
      (src034[42] << 34) +
      (src034[43] << 34) +
      (src034[44] << 34) +
      (src034[45] << 34) +
      (src034[46] << 34) +
      (src034[47] << 34) +
      (src034[48] << 34) +
      (src034[49] << 34) +
      (src034[50] << 34) +
      (src034[51] << 34) +
      (src034[52] << 34) +
      (src034[53] << 34) +
      (src034[54] << 34) +
      (src034[55] << 34) +
      (src034[56] << 34) +
      (src034[57] << 34) +
      (src034[58] << 34) +
      (src034[59] << 34) +
      (src034[60] << 34) +
      (src034[61] << 34) +
      (src034[62] << 34) +
      (src034[63] << 34) +
      (src034[64] << 34) +
      (src034[65] << 34) +
      (src034[66] << 34) +
      (src034[67] << 34) +
      (src034[68] << 34) +
      (src034[69] << 34) +
      (src034[70] << 34) +
      (src034[71] << 34) +
      (src034[72] << 34) +
      (src034[73] << 34) +
      (src034[74] << 34) +
      (src034[75] << 34) +
      (src034[76] << 34) +
      (src034[77] << 34) +
      (src034[78] << 34) +
      (src034[79] << 34) +
      (src034[80] << 34) +
      (src034[81] << 34) +
      (src034[82] << 34) +
      (src034[83] << 34) +
      (src034[84] << 34) +
      (src034[85] << 34) +
      (src034[86] << 34) +
      (src034[87] << 34) +
      (src034[88] << 34) +
      (src034[89] << 34) +
      (src034[90] << 34) +
      (src034[91] << 34) +
      (src034[92] << 34) +
      (src034[93] << 34) +
      (src034[94] << 34) +
      (src034[95] << 34) +
      (src034[96] << 34) +
      (src034[97] << 34) +
      (src034[98] << 34) +
      (src034[99] << 34) +
      (src034[100] << 34) +
      (src034[101] << 34) +
      (src034[102] << 34) +
      (src034[103] << 34) +
      (src034[104] << 34) +
      (src034[105] << 34) +
      (src034[106] << 34) +
      (src034[107] << 34) +
      (src034[108] << 34) +
      (src034[109] << 34) +
      (src034[110] << 34) +
      (src034[111] << 34) +
      (src034[112] << 34) +
      (src034[113] << 34) +
      (src034[114] << 34) +
      (src034[115] << 34) +
      (src034[116] << 34) +
      (src034[117] << 34) +
      (src034[118] << 34) +
      (src034[119] << 34) +
      (src034[120] << 34) +
      (src034[121] << 34) +
      (src034[122] << 34) +
      (src034[123] << 34) +
      (src034[124] << 34) +
      (src034[125] << 34) +
      (src034[126] << 34) +
      (src034[127] << 34) +
      (src035[0] << 35) +
      (src035[1] << 35) +
      (src035[2] << 35) +
      (src035[3] << 35) +
      (src035[4] << 35) +
      (src035[5] << 35) +
      (src035[6] << 35) +
      (src035[7] << 35) +
      (src035[8] << 35) +
      (src035[9] << 35) +
      (src035[10] << 35) +
      (src035[11] << 35) +
      (src035[12] << 35) +
      (src035[13] << 35) +
      (src035[14] << 35) +
      (src035[15] << 35) +
      (src035[16] << 35) +
      (src035[17] << 35) +
      (src035[18] << 35) +
      (src035[19] << 35) +
      (src035[20] << 35) +
      (src035[21] << 35) +
      (src035[22] << 35) +
      (src035[23] << 35) +
      (src035[24] << 35) +
      (src035[25] << 35) +
      (src035[26] << 35) +
      (src035[27] << 35) +
      (src035[28] << 35) +
      (src035[29] << 35) +
      (src035[30] << 35) +
      (src035[31] << 35) +
      (src035[32] << 35) +
      (src035[33] << 35) +
      (src035[34] << 35) +
      (src035[35] << 35) +
      (src035[36] << 35) +
      (src035[37] << 35) +
      (src035[38] << 35) +
      (src035[39] << 35) +
      (src035[40] << 35) +
      (src035[41] << 35) +
      (src035[42] << 35) +
      (src035[43] << 35) +
      (src035[44] << 35) +
      (src035[45] << 35) +
      (src035[46] << 35) +
      (src035[47] << 35) +
      (src035[48] << 35) +
      (src035[49] << 35) +
      (src035[50] << 35) +
      (src035[51] << 35) +
      (src035[52] << 35) +
      (src035[53] << 35) +
      (src035[54] << 35) +
      (src035[55] << 35) +
      (src035[56] << 35) +
      (src035[57] << 35) +
      (src035[58] << 35) +
      (src035[59] << 35) +
      (src035[60] << 35) +
      (src035[61] << 35) +
      (src035[62] << 35) +
      (src035[63] << 35) +
      (src035[64] << 35) +
      (src035[65] << 35) +
      (src035[66] << 35) +
      (src035[67] << 35) +
      (src035[68] << 35) +
      (src035[69] << 35) +
      (src035[70] << 35) +
      (src035[71] << 35) +
      (src035[72] << 35) +
      (src035[73] << 35) +
      (src035[74] << 35) +
      (src035[75] << 35) +
      (src035[76] << 35) +
      (src035[77] << 35) +
      (src035[78] << 35) +
      (src035[79] << 35) +
      (src035[80] << 35) +
      (src035[81] << 35) +
      (src035[82] << 35) +
      (src035[83] << 35) +
      (src035[84] << 35) +
      (src035[85] << 35) +
      (src035[86] << 35) +
      (src035[87] << 35) +
      (src035[88] << 35) +
      (src035[89] << 35) +
      (src035[90] << 35) +
      (src035[91] << 35) +
      (src035[92] << 35) +
      (src035[93] << 35) +
      (src035[94] << 35) +
      (src035[95] << 35) +
      (src035[96] << 35) +
      (src035[97] << 35) +
      (src035[98] << 35) +
      (src035[99] << 35) +
      (src035[100] << 35) +
      (src035[101] << 35) +
      (src035[102] << 35) +
      (src035[103] << 35) +
      (src035[104] << 35) +
      (src035[105] << 35) +
      (src035[106] << 35) +
      (src035[107] << 35) +
      (src035[108] << 35) +
      (src035[109] << 35) +
      (src035[110] << 35) +
      (src035[111] << 35) +
      (src035[112] << 35) +
      (src035[113] << 35) +
      (src035[114] << 35) +
      (src035[115] << 35) +
      (src035[116] << 35) +
      (src035[117] << 35) +
      (src035[118] << 35) +
      (src035[119] << 35) +
      (src035[120] << 35) +
      (src035[121] << 35) +
      (src035[122] << 35) +
      (src035[123] << 35) +
      (src035[124] << 35) +
      (src035[125] << 35) +
      (src035[126] << 35) +
      (src035[127] << 35) +
      (src036[0] << 36) +
      (src036[1] << 36) +
      (src036[2] << 36) +
      (src036[3] << 36) +
      (src036[4] << 36) +
      (src036[5] << 36) +
      (src036[6] << 36) +
      (src036[7] << 36) +
      (src036[8] << 36) +
      (src036[9] << 36) +
      (src036[10] << 36) +
      (src036[11] << 36) +
      (src036[12] << 36) +
      (src036[13] << 36) +
      (src036[14] << 36) +
      (src036[15] << 36) +
      (src036[16] << 36) +
      (src036[17] << 36) +
      (src036[18] << 36) +
      (src036[19] << 36) +
      (src036[20] << 36) +
      (src036[21] << 36) +
      (src036[22] << 36) +
      (src036[23] << 36) +
      (src036[24] << 36) +
      (src036[25] << 36) +
      (src036[26] << 36) +
      (src036[27] << 36) +
      (src036[28] << 36) +
      (src036[29] << 36) +
      (src036[30] << 36) +
      (src036[31] << 36) +
      (src036[32] << 36) +
      (src036[33] << 36) +
      (src036[34] << 36) +
      (src036[35] << 36) +
      (src036[36] << 36) +
      (src036[37] << 36) +
      (src036[38] << 36) +
      (src036[39] << 36) +
      (src036[40] << 36) +
      (src036[41] << 36) +
      (src036[42] << 36) +
      (src036[43] << 36) +
      (src036[44] << 36) +
      (src036[45] << 36) +
      (src036[46] << 36) +
      (src036[47] << 36) +
      (src036[48] << 36) +
      (src036[49] << 36) +
      (src036[50] << 36) +
      (src036[51] << 36) +
      (src036[52] << 36) +
      (src036[53] << 36) +
      (src036[54] << 36) +
      (src036[55] << 36) +
      (src036[56] << 36) +
      (src036[57] << 36) +
      (src036[58] << 36) +
      (src036[59] << 36) +
      (src036[60] << 36) +
      (src036[61] << 36) +
      (src036[62] << 36) +
      (src036[63] << 36) +
      (src036[64] << 36) +
      (src036[65] << 36) +
      (src036[66] << 36) +
      (src036[67] << 36) +
      (src036[68] << 36) +
      (src036[69] << 36) +
      (src036[70] << 36) +
      (src036[71] << 36) +
      (src036[72] << 36) +
      (src036[73] << 36) +
      (src036[74] << 36) +
      (src036[75] << 36) +
      (src036[76] << 36) +
      (src036[77] << 36) +
      (src036[78] << 36) +
      (src036[79] << 36) +
      (src036[80] << 36) +
      (src036[81] << 36) +
      (src036[82] << 36) +
      (src036[83] << 36) +
      (src036[84] << 36) +
      (src036[85] << 36) +
      (src036[86] << 36) +
      (src036[87] << 36) +
      (src036[88] << 36) +
      (src036[89] << 36) +
      (src036[90] << 36) +
      (src036[91] << 36) +
      (src036[92] << 36) +
      (src036[93] << 36) +
      (src036[94] << 36) +
      (src036[95] << 36) +
      (src036[96] << 36) +
      (src036[97] << 36) +
      (src036[98] << 36) +
      (src036[99] << 36) +
      (src036[100] << 36) +
      (src036[101] << 36) +
      (src036[102] << 36) +
      (src036[103] << 36) +
      (src036[104] << 36) +
      (src036[105] << 36) +
      (src036[106] << 36) +
      (src036[107] << 36) +
      (src036[108] << 36) +
      (src036[109] << 36) +
      (src036[110] << 36) +
      (src036[111] << 36) +
      (src036[112] << 36) +
      (src036[113] << 36) +
      (src036[114] << 36) +
      (src036[115] << 36) +
      (src036[116] << 36) +
      (src036[117] << 36) +
      (src036[118] << 36) +
      (src036[119] << 36) +
      (src036[120] << 36) +
      (src036[121] << 36) +
      (src036[122] << 36) +
      (src036[123] << 36) +
      (src036[124] << 36) +
      (src036[125] << 36) +
      (src036[126] << 36) +
      (src036[127] << 36) +
      (src037[0] << 37) +
      (src037[1] << 37) +
      (src037[2] << 37) +
      (src037[3] << 37) +
      (src037[4] << 37) +
      (src037[5] << 37) +
      (src037[6] << 37) +
      (src037[7] << 37) +
      (src037[8] << 37) +
      (src037[9] << 37) +
      (src037[10] << 37) +
      (src037[11] << 37) +
      (src037[12] << 37) +
      (src037[13] << 37) +
      (src037[14] << 37) +
      (src037[15] << 37) +
      (src037[16] << 37) +
      (src037[17] << 37) +
      (src037[18] << 37) +
      (src037[19] << 37) +
      (src037[20] << 37) +
      (src037[21] << 37) +
      (src037[22] << 37) +
      (src037[23] << 37) +
      (src037[24] << 37) +
      (src037[25] << 37) +
      (src037[26] << 37) +
      (src037[27] << 37) +
      (src037[28] << 37) +
      (src037[29] << 37) +
      (src037[30] << 37) +
      (src037[31] << 37) +
      (src037[32] << 37) +
      (src037[33] << 37) +
      (src037[34] << 37) +
      (src037[35] << 37) +
      (src037[36] << 37) +
      (src037[37] << 37) +
      (src037[38] << 37) +
      (src037[39] << 37) +
      (src037[40] << 37) +
      (src037[41] << 37) +
      (src037[42] << 37) +
      (src037[43] << 37) +
      (src037[44] << 37) +
      (src037[45] << 37) +
      (src037[46] << 37) +
      (src037[47] << 37) +
      (src037[48] << 37) +
      (src037[49] << 37) +
      (src037[50] << 37) +
      (src037[51] << 37) +
      (src037[52] << 37) +
      (src037[53] << 37) +
      (src037[54] << 37) +
      (src037[55] << 37) +
      (src037[56] << 37) +
      (src037[57] << 37) +
      (src037[58] << 37) +
      (src037[59] << 37) +
      (src037[60] << 37) +
      (src037[61] << 37) +
      (src037[62] << 37) +
      (src037[63] << 37) +
      (src037[64] << 37) +
      (src037[65] << 37) +
      (src037[66] << 37) +
      (src037[67] << 37) +
      (src037[68] << 37) +
      (src037[69] << 37) +
      (src037[70] << 37) +
      (src037[71] << 37) +
      (src037[72] << 37) +
      (src037[73] << 37) +
      (src037[74] << 37) +
      (src037[75] << 37) +
      (src037[76] << 37) +
      (src037[77] << 37) +
      (src037[78] << 37) +
      (src037[79] << 37) +
      (src037[80] << 37) +
      (src037[81] << 37) +
      (src037[82] << 37) +
      (src037[83] << 37) +
      (src037[84] << 37) +
      (src037[85] << 37) +
      (src037[86] << 37) +
      (src037[87] << 37) +
      (src037[88] << 37) +
      (src037[89] << 37) +
      (src037[90] << 37) +
      (src037[91] << 37) +
      (src037[92] << 37) +
      (src037[93] << 37) +
      (src037[94] << 37) +
      (src037[95] << 37) +
      (src037[96] << 37) +
      (src037[97] << 37) +
      (src037[98] << 37) +
      (src037[99] << 37) +
      (src037[100] << 37) +
      (src037[101] << 37) +
      (src037[102] << 37) +
      (src037[103] << 37) +
      (src037[104] << 37) +
      (src037[105] << 37) +
      (src037[106] << 37) +
      (src037[107] << 37) +
      (src037[108] << 37) +
      (src037[109] << 37) +
      (src037[110] << 37) +
      (src037[111] << 37) +
      (src037[112] << 37) +
      (src037[113] << 37) +
      (src037[114] << 37) +
      (src037[115] << 37) +
      (src037[116] << 37) +
      (src037[117] << 37) +
      (src037[118] << 37) +
      (src037[119] << 37) +
      (src037[120] << 37) +
      (src037[121] << 37) +
      (src037[122] << 37) +
      (src037[123] << 37) +
      (src037[124] << 37) +
      (src037[125] << 37) +
      (src037[126] << 37) +
      (src037[127] << 37) +
      (src038[0] << 38) +
      (src038[1] << 38) +
      (src038[2] << 38) +
      (src038[3] << 38) +
      (src038[4] << 38) +
      (src038[5] << 38) +
      (src038[6] << 38) +
      (src038[7] << 38) +
      (src038[8] << 38) +
      (src038[9] << 38) +
      (src038[10] << 38) +
      (src038[11] << 38) +
      (src038[12] << 38) +
      (src038[13] << 38) +
      (src038[14] << 38) +
      (src038[15] << 38) +
      (src038[16] << 38) +
      (src038[17] << 38) +
      (src038[18] << 38) +
      (src038[19] << 38) +
      (src038[20] << 38) +
      (src038[21] << 38) +
      (src038[22] << 38) +
      (src038[23] << 38) +
      (src038[24] << 38) +
      (src038[25] << 38) +
      (src038[26] << 38) +
      (src038[27] << 38) +
      (src038[28] << 38) +
      (src038[29] << 38) +
      (src038[30] << 38) +
      (src038[31] << 38) +
      (src038[32] << 38) +
      (src038[33] << 38) +
      (src038[34] << 38) +
      (src038[35] << 38) +
      (src038[36] << 38) +
      (src038[37] << 38) +
      (src038[38] << 38) +
      (src038[39] << 38) +
      (src038[40] << 38) +
      (src038[41] << 38) +
      (src038[42] << 38) +
      (src038[43] << 38) +
      (src038[44] << 38) +
      (src038[45] << 38) +
      (src038[46] << 38) +
      (src038[47] << 38) +
      (src038[48] << 38) +
      (src038[49] << 38) +
      (src038[50] << 38) +
      (src038[51] << 38) +
      (src038[52] << 38) +
      (src038[53] << 38) +
      (src038[54] << 38) +
      (src038[55] << 38) +
      (src038[56] << 38) +
      (src038[57] << 38) +
      (src038[58] << 38) +
      (src038[59] << 38) +
      (src038[60] << 38) +
      (src038[61] << 38) +
      (src038[62] << 38) +
      (src038[63] << 38) +
      (src038[64] << 38) +
      (src038[65] << 38) +
      (src038[66] << 38) +
      (src038[67] << 38) +
      (src038[68] << 38) +
      (src038[69] << 38) +
      (src038[70] << 38) +
      (src038[71] << 38) +
      (src038[72] << 38) +
      (src038[73] << 38) +
      (src038[74] << 38) +
      (src038[75] << 38) +
      (src038[76] << 38) +
      (src038[77] << 38) +
      (src038[78] << 38) +
      (src038[79] << 38) +
      (src038[80] << 38) +
      (src038[81] << 38) +
      (src038[82] << 38) +
      (src038[83] << 38) +
      (src038[84] << 38) +
      (src038[85] << 38) +
      (src038[86] << 38) +
      (src038[87] << 38) +
      (src038[88] << 38) +
      (src038[89] << 38) +
      (src038[90] << 38) +
      (src038[91] << 38) +
      (src038[92] << 38) +
      (src038[93] << 38) +
      (src038[94] << 38) +
      (src038[95] << 38) +
      (src038[96] << 38) +
      (src038[97] << 38) +
      (src038[98] << 38) +
      (src038[99] << 38) +
      (src038[100] << 38) +
      (src038[101] << 38) +
      (src038[102] << 38) +
      (src038[103] << 38) +
      (src038[104] << 38) +
      (src038[105] << 38) +
      (src038[106] << 38) +
      (src038[107] << 38) +
      (src038[108] << 38) +
      (src038[109] << 38) +
      (src038[110] << 38) +
      (src038[111] << 38) +
      (src038[112] << 38) +
      (src038[113] << 38) +
      (src038[114] << 38) +
      (src038[115] << 38) +
      (src038[116] << 38) +
      (src038[117] << 38) +
      (src038[118] << 38) +
      (src038[119] << 38) +
      (src038[120] << 38) +
      (src038[121] << 38) +
      (src038[122] << 38) +
      (src038[123] << 38) +
      (src038[124] << 38) +
      (src038[125] << 38) +
      (src038[126] << 38) +
      (src038[127] << 38) +
      (src039[0] << 39) +
      (src039[1] << 39) +
      (src039[2] << 39) +
      (src039[3] << 39) +
      (src039[4] << 39) +
      (src039[5] << 39) +
      (src039[6] << 39) +
      (src039[7] << 39) +
      (src039[8] << 39) +
      (src039[9] << 39) +
      (src039[10] << 39) +
      (src039[11] << 39) +
      (src039[12] << 39) +
      (src039[13] << 39) +
      (src039[14] << 39) +
      (src039[15] << 39) +
      (src039[16] << 39) +
      (src039[17] << 39) +
      (src039[18] << 39) +
      (src039[19] << 39) +
      (src039[20] << 39) +
      (src039[21] << 39) +
      (src039[22] << 39) +
      (src039[23] << 39) +
      (src039[24] << 39) +
      (src039[25] << 39) +
      (src039[26] << 39) +
      (src039[27] << 39) +
      (src039[28] << 39) +
      (src039[29] << 39) +
      (src039[30] << 39) +
      (src039[31] << 39) +
      (src039[32] << 39) +
      (src039[33] << 39) +
      (src039[34] << 39) +
      (src039[35] << 39) +
      (src039[36] << 39) +
      (src039[37] << 39) +
      (src039[38] << 39) +
      (src039[39] << 39) +
      (src039[40] << 39) +
      (src039[41] << 39) +
      (src039[42] << 39) +
      (src039[43] << 39) +
      (src039[44] << 39) +
      (src039[45] << 39) +
      (src039[46] << 39) +
      (src039[47] << 39) +
      (src039[48] << 39) +
      (src039[49] << 39) +
      (src039[50] << 39) +
      (src039[51] << 39) +
      (src039[52] << 39) +
      (src039[53] << 39) +
      (src039[54] << 39) +
      (src039[55] << 39) +
      (src039[56] << 39) +
      (src039[57] << 39) +
      (src039[58] << 39) +
      (src039[59] << 39) +
      (src039[60] << 39) +
      (src039[61] << 39) +
      (src039[62] << 39) +
      (src039[63] << 39) +
      (src039[64] << 39) +
      (src039[65] << 39) +
      (src039[66] << 39) +
      (src039[67] << 39) +
      (src039[68] << 39) +
      (src039[69] << 39) +
      (src039[70] << 39) +
      (src039[71] << 39) +
      (src039[72] << 39) +
      (src039[73] << 39) +
      (src039[74] << 39) +
      (src039[75] << 39) +
      (src039[76] << 39) +
      (src039[77] << 39) +
      (src039[78] << 39) +
      (src039[79] << 39) +
      (src039[80] << 39) +
      (src039[81] << 39) +
      (src039[82] << 39) +
      (src039[83] << 39) +
      (src039[84] << 39) +
      (src039[85] << 39) +
      (src039[86] << 39) +
      (src039[87] << 39) +
      (src039[88] << 39) +
      (src039[89] << 39) +
      (src039[90] << 39) +
      (src039[91] << 39) +
      (src039[92] << 39) +
      (src039[93] << 39) +
      (src039[94] << 39) +
      (src039[95] << 39) +
      (src039[96] << 39) +
      (src039[97] << 39) +
      (src039[98] << 39) +
      (src039[99] << 39) +
      (src039[100] << 39) +
      (src039[101] << 39) +
      (src039[102] << 39) +
      (src039[103] << 39) +
      (src039[104] << 39) +
      (src039[105] << 39) +
      (src039[106] << 39) +
      (src039[107] << 39) +
      (src039[108] << 39) +
      (src039[109] << 39) +
      (src039[110] << 39) +
      (src039[111] << 39) +
      (src039[112] << 39) +
      (src039[113] << 39) +
      (src039[114] << 39) +
      (src039[115] << 39) +
      (src039[116] << 39) +
      (src039[117] << 39) +
      (src039[118] << 39) +
      (src039[119] << 39) +
      (src039[120] << 39) +
      (src039[121] << 39) +
      (src039[122] << 39) +
      (src039[123] << 39) +
      (src039[124] << 39) +
      (src039[125] << 39) +
      (src039[126] << 39) +
      (src039[127] << 39) +
      (src040[0] << 40) +
      (src040[1] << 40) +
      (src040[2] << 40) +
      (src040[3] << 40) +
      (src040[4] << 40) +
      (src040[5] << 40) +
      (src040[6] << 40) +
      (src040[7] << 40) +
      (src040[8] << 40) +
      (src040[9] << 40) +
      (src040[10] << 40) +
      (src040[11] << 40) +
      (src040[12] << 40) +
      (src040[13] << 40) +
      (src040[14] << 40) +
      (src040[15] << 40) +
      (src040[16] << 40) +
      (src040[17] << 40) +
      (src040[18] << 40) +
      (src040[19] << 40) +
      (src040[20] << 40) +
      (src040[21] << 40) +
      (src040[22] << 40) +
      (src040[23] << 40) +
      (src040[24] << 40) +
      (src040[25] << 40) +
      (src040[26] << 40) +
      (src040[27] << 40) +
      (src040[28] << 40) +
      (src040[29] << 40) +
      (src040[30] << 40) +
      (src040[31] << 40) +
      (src040[32] << 40) +
      (src040[33] << 40) +
      (src040[34] << 40) +
      (src040[35] << 40) +
      (src040[36] << 40) +
      (src040[37] << 40) +
      (src040[38] << 40) +
      (src040[39] << 40) +
      (src040[40] << 40) +
      (src040[41] << 40) +
      (src040[42] << 40) +
      (src040[43] << 40) +
      (src040[44] << 40) +
      (src040[45] << 40) +
      (src040[46] << 40) +
      (src040[47] << 40) +
      (src040[48] << 40) +
      (src040[49] << 40) +
      (src040[50] << 40) +
      (src040[51] << 40) +
      (src040[52] << 40) +
      (src040[53] << 40) +
      (src040[54] << 40) +
      (src040[55] << 40) +
      (src040[56] << 40) +
      (src040[57] << 40) +
      (src040[58] << 40) +
      (src040[59] << 40) +
      (src040[60] << 40) +
      (src040[61] << 40) +
      (src040[62] << 40) +
      (src040[63] << 40) +
      (src040[64] << 40) +
      (src040[65] << 40) +
      (src040[66] << 40) +
      (src040[67] << 40) +
      (src040[68] << 40) +
      (src040[69] << 40) +
      (src040[70] << 40) +
      (src040[71] << 40) +
      (src040[72] << 40) +
      (src040[73] << 40) +
      (src040[74] << 40) +
      (src040[75] << 40) +
      (src040[76] << 40) +
      (src040[77] << 40) +
      (src040[78] << 40) +
      (src040[79] << 40) +
      (src040[80] << 40) +
      (src040[81] << 40) +
      (src040[82] << 40) +
      (src040[83] << 40) +
      (src040[84] << 40) +
      (src040[85] << 40) +
      (src040[86] << 40) +
      (src040[87] << 40) +
      (src040[88] << 40) +
      (src040[89] << 40) +
      (src040[90] << 40) +
      (src040[91] << 40) +
      (src040[92] << 40) +
      (src040[93] << 40) +
      (src040[94] << 40) +
      (src040[95] << 40) +
      (src040[96] << 40) +
      (src040[97] << 40) +
      (src040[98] << 40) +
      (src040[99] << 40) +
      (src040[100] << 40) +
      (src040[101] << 40) +
      (src040[102] << 40) +
      (src040[103] << 40) +
      (src040[104] << 40) +
      (src040[105] << 40) +
      (src040[106] << 40) +
      (src040[107] << 40) +
      (src040[108] << 40) +
      (src040[109] << 40) +
      (src040[110] << 40) +
      (src040[111] << 40) +
      (src040[112] << 40) +
      (src040[113] << 40) +
      (src040[114] << 40) +
      (src040[115] << 40) +
      (src040[116] << 40) +
      (src040[117] << 40) +
      (src040[118] << 40) +
      (src040[119] << 40) +
      (src040[120] << 40) +
      (src040[121] << 40) +
      (src040[122] << 40) +
      (src040[123] << 40) +
      (src040[124] << 40) +
      (src040[125] << 40) +
      (src040[126] << 40) +
      (src040[127] << 40) +
      (src041[0] << 41) +
      (src041[1] << 41) +
      (src041[2] << 41) +
      (src041[3] << 41) +
      (src041[4] << 41) +
      (src041[5] << 41) +
      (src041[6] << 41) +
      (src041[7] << 41) +
      (src041[8] << 41) +
      (src041[9] << 41) +
      (src041[10] << 41) +
      (src041[11] << 41) +
      (src041[12] << 41) +
      (src041[13] << 41) +
      (src041[14] << 41) +
      (src041[15] << 41) +
      (src041[16] << 41) +
      (src041[17] << 41) +
      (src041[18] << 41) +
      (src041[19] << 41) +
      (src041[20] << 41) +
      (src041[21] << 41) +
      (src041[22] << 41) +
      (src041[23] << 41) +
      (src041[24] << 41) +
      (src041[25] << 41) +
      (src041[26] << 41) +
      (src041[27] << 41) +
      (src041[28] << 41) +
      (src041[29] << 41) +
      (src041[30] << 41) +
      (src041[31] << 41) +
      (src041[32] << 41) +
      (src041[33] << 41) +
      (src041[34] << 41) +
      (src041[35] << 41) +
      (src041[36] << 41) +
      (src041[37] << 41) +
      (src041[38] << 41) +
      (src041[39] << 41) +
      (src041[40] << 41) +
      (src041[41] << 41) +
      (src041[42] << 41) +
      (src041[43] << 41) +
      (src041[44] << 41) +
      (src041[45] << 41) +
      (src041[46] << 41) +
      (src041[47] << 41) +
      (src041[48] << 41) +
      (src041[49] << 41) +
      (src041[50] << 41) +
      (src041[51] << 41) +
      (src041[52] << 41) +
      (src041[53] << 41) +
      (src041[54] << 41) +
      (src041[55] << 41) +
      (src041[56] << 41) +
      (src041[57] << 41) +
      (src041[58] << 41) +
      (src041[59] << 41) +
      (src041[60] << 41) +
      (src041[61] << 41) +
      (src041[62] << 41) +
      (src041[63] << 41) +
      (src041[64] << 41) +
      (src041[65] << 41) +
      (src041[66] << 41) +
      (src041[67] << 41) +
      (src041[68] << 41) +
      (src041[69] << 41) +
      (src041[70] << 41) +
      (src041[71] << 41) +
      (src041[72] << 41) +
      (src041[73] << 41) +
      (src041[74] << 41) +
      (src041[75] << 41) +
      (src041[76] << 41) +
      (src041[77] << 41) +
      (src041[78] << 41) +
      (src041[79] << 41) +
      (src041[80] << 41) +
      (src041[81] << 41) +
      (src041[82] << 41) +
      (src041[83] << 41) +
      (src041[84] << 41) +
      (src041[85] << 41) +
      (src041[86] << 41) +
      (src041[87] << 41) +
      (src041[88] << 41) +
      (src041[89] << 41) +
      (src041[90] << 41) +
      (src041[91] << 41) +
      (src041[92] << 41) +
      (src041[93] << 41) +
      (src041[94] << 41) +
      (src041[95] << 41) +
      (src041[96] << 41) +
      (src041[97] << 41) +
      (src041[98] << 41) +
      (src041[99] << 41) +
      (src041[100] << 41) +
      (src041[101] << 41) +
      (src041[102] << 41) +
      (src041[103] << 41) +
      (src041[104] << 41) +
      (src041[105] << 41) +
      (src041[106] << 41) +
      (src041[107] << 41) +
      (src041[108] << 41) +
      (src041[109] << 41) +
      (src041[110] << 41) +
      (src041[111] << 41) +
      (src041[112] << 41) +
      (src041[113] << 41) +
      (src041[114] << 41) +
      (src041[115] << 41) +
      (src041[116] << 41) +
      (src041[117] << 41) +
      (src041[118] << 41) +
      (src041[119] << 41) +
      (src041[120] << 41) +
      (src041[121] << 41) +
      (src041[122] << 41) +
      (src041[123] << 41) +
      (src041[124] << 41) +
      (src041[125] << 41) +
      (src041[126] << 41) +
      (src041[127] << 41) +
      (src042[0] << 42) +
      (src042[1] << 42) +
      (src042[2] << 42) +
      (src042[3] << 42) +
      (src042[4] << 42) +
      (src042[5] << 42) +
      (src042[6] << 42) +
      (src042[7] << 42) +
      (src042[8] << 42) +
      (src042[9] << 42) +
      (src042[10] << 42) +
      (src042[11] << 42) +
      (src042[12] << 42) +
      (src042[13] << 42) +
      (src042[14] << 42) +
      (src042[15] << 42) +
      (src042[16] << 42) +
      (src042[17] << 42) +
      (src042[18] << 42) +
      (src042[19] << 42) +
      (src042[20] << 42) +
      (src042[21] << 42) +
      (src042[22] << 42) +
      (src042[23] << 42) +
      (src042[24] << 42) +
      (src042[25] << 42) +
      (src042[26] << 42) +
      (src042[27] << 42) +
      (src042[28] << 42) +
      (src042[29] << 42) +
      (src042[30] << 42) +
      (src042[31] << 42) +
      (src042[32] << 42) +
      (src042[33] << 42) +
      (src042[34] << 42) +
      (src042[35] << 42) +
      (src042[36] << 42) +
      (src042[37] << 42) +
      (src042[38] << 42) +
      (src042[39] << 42) +
      (src042[40] << 42) +
      (src042[41] << 42) +
      (src042[42] << 42) +
      (src042[43] << 42) +
      (src042[44] << 42) +
      (src042[45] << 42) +
      (src042[46] << 42) +
      (src042[47] << 42) +
      (src042[48] << 42) +
      (src042[49] << 42) +
      (src042[50] << 42) +
      (src042[51] << 42) +
      (src042[52] << 42) +
      (src042[53] << 42) +
      (src042[54] << 42) +
      (src042[55] << 42) +
      (src042[56] << 42) +
      (src042[57] << 42) +
      (src042[58] << 42) +
      (src042[59] << 42) +
      (src042[60] << 42) +
      (src042[61] << 42) +
      (src042[62] << 42) +
      (src042[63] << 42) +
      (src042[64] << 42) +
      (src042[65] << 42) +
      (src042[66] << 42) +
      (src042[67] << 42) +
      (src042[68] << 42) +
      (src042[69] << 42) +
      (src042[70] << 42) +
      (src042[71] << 42) +
      (src042[72] << 42) +
      (src042[73] << 42) +
      (src042[74] << 42) +
      (src042[75] << 42) +
      (src042[76] << 42) +
      (src042[77] << 42) +
      (src042[78] << 42) +
      (src042[79] << 42) +
      (src042[80] << 42) +
      (src042[81] << 42) +
      (src042[82] << 42) +
      (src042[83] << 42) +
      (src042[84] << 42) +
      (src042[85] << 42) +
      (src042[86] << 42) +
      (src042[87] << 42) +
      (src042[88] << 42) +
      (src042[89] << 42) +
      (src042[90] << 42) +
      (src042[91] << 42) +
      (src042[92] << 42) +
      (src042[93] << 42) +
      (src042[94] << 42) +
      (src042[95] << 42) +
      (src042[96] << 42) +
      (src042[97] << 42) +
      (src042[98] << 42) +
      (src042[99] << 42) +
      (src042[100] << 42) +
      (src042[101] << 42) +
      (src042[102] << 42) +
      (src042[103] << 42) +
      (src042[104] << 42) +
      (src042[105] << 42) +
      (src042[106] << 42) +
      (src042[107] << 42) +
      (src042[108] << 42) +
      (src042[109] << 42) +
      (src042[110] << 42) +
      (src042[111] << 42) +
      (src042[112] << 42) +
      (src042[113] << 42) +
      (src042[114] << 42) +
      (src042[115] << 42) +
      (src042[116] << 42) +
      (src042[117] << 42) +
      (src042[118] << 42) +
      (src042[119] << 42) +
      (src042[120] << 42) +
      (src042[121] << 42) +
      (src042[122] << 42) +
      (src042[123] << 42) +
      (src042[124] << 42) +
      (src042[125] << 42) +
      (src042[126] << 42) +
      (src042[127] << 42) +
      (src043[0] << 43) +
      (src043[1] << 43) +
      (src043[2] << 43) +
      (src043[3] << 43) +
      (src043[4] << 43) +
      (src043[5] << 43) +
      (src043[6] << 43) +
      (src043[7] << 43) +
      (src043[8] << 43) +
      (src043[9] << 43) +
      (src043[10] << 43) +
      (src043[11] << 43) +
      (src043[12] << 43) +
      (src043[13] << 43) +
      (src043[14] << 43) +
      (src043[15] << 43) +
      (src043[16] << 43) +
      (src043[17] << 43) +
      (src043[18] << 43) +
      (src043[19] << 43) +
      (src043[20] << 43) +
      (src043[21] << 43) +
      (src043[22] << 43) +
      (src043[23] << 43) +
      (src043[24] << 43) +
      (src043[25] << 43) +
      (src043[26] << 43) +
      (src043[27] << 43) +
      (src043[28] << 43) +
      (src043[29] << 43) +
      (src043[30] << 43) +
      (src043[31] << 43) +
      (src043[32] << 43) +
      (src043[33] << 43) +
      (src043[34] << 43) +
      (src043[35] << 43) +
      (src043[36] << 43) +
      (src043[37] << 43) +
      (src043[38] << 43) +
      (src043[39] << 43) +
      (src043[40] << 43) +
      (src043[41] << 43) +
      (src043[42] << 43) +
      (src043[43] << 43) +
      (src043[44] << 43) +
      (src043[45] << 43) +
      (src043[46] << 43) +
      (src043[47] << 43) +
      (src043[48] << 43) +
      (src043[49] << 43) +
      (src043[50] << 43) +
      (src043[51] << 43) +
      (src043[52] << 43) +
      (src043[53] << 43) +
      (src043[54] << 43) +
      (src043[55] << 43) +
      (src043[56] << 43) +
      (src043[57] << 43) +
      (src043[58] << 43) +
      (src043[59] << 43) +
      (src043[60] << 43) +
      (src043[61] << 43) +
      (src043[62] << 43) +
      (src043[63] << 43) +
      (src043[64] << 43) +
      (src043[65] << 43) +
      (src043[66] << 43) +
      (src043[67] << 43) +
      (src043[68] << 43) +
      (src043[69] << 43) +
      (src043[70] << 43) +
      (src043[71] << 43) +
      (src043[72] << 43) +
      (src043[73] << 43) +
      (src043[74] << 43) +
      (src043[75] << 43) +
      (src043[76] << 43) +
      (src043[77] << 43) +
      (src043[78] << 43) +
      (src043[79] << 43) +
      (src043[80] << 43) +
      (src043[81] << 43) +
      (src043[82] << 43) +
      (src043[83] << 43) +
      (src043[84] << 43) +
      (src043[85] << 43) +
      (src043[86] << 43) +
      (src043[87] << 43) +
      (src043[88] << 43) +
      (src043[89] << 43) +
      (src043[90] << 43) +
      (src043[91] << 43) +
      (src043[92] << 43) +
      (src043[93] << 43) +
      (src043[94] << 43) +
      (src043[95] << 43) +
      (src043[96] << 43) +
      (src043[97] << 43) +
      (src043[98] << 43) +
      (src043[99] << 43) +
      (src043[100] << 43) +
      (src043[101] << 43) +
      (src043[102] << 43) +
      (src043[103] << 43) +
      (src043[104] << 43) +
      (src043[105] << 43) +
      (src043[106] << 43) +
      (src043[107] << 43) +
      (src043[108] << 43) +
      (src043[109] << 43) +
      (src043[110] << 43) +
      (src043[111] << 43) +
      (src043[112] << 43) +
      (src043[113] << 43) +
      (src043[114] << 43) +
      (src043[115] << 43) +
      (src043[116] << 43) +
      (src043[117] << 43) +
      (src043[118] << 43) +
      (src043[119] << 43) +
      (src043[120] << 43) +
      (src043[121] << 43) +
      (src043[122] << 43) +
      (src043[123] << 43) +
      (src043[124] << 43) +
      (src043[125] << 43) +
      (src043[126] << 43) +
      (src043[127] << 43) +
      (src044[0] << 44) +
      (src044[1] << 44) +
      (src044[2] << 44) +
      (src044[3] << 44) +
      (src044[4] << 44) +
      (src044[5] << 44) +
      (src044[6] << 44) +
      (src044[7] << 44) +
      (src044[8] << 44) +
      (src044[9] << 44) +
      (src044[10] << 44) +
      (src044[11] << 44) +
      (src044[12] << 44) +
      (src044[13] << 44) +
      (src044[14] << 44) +
      (src044[15] << 44) +
      (src044[16] << 44) +
      (src044[17] << 44) +
      (src044[18] << 44) +
      (src044[19] << 44) +
      (src044[20] << 44) +
      (src044[21] << 44) +
      (src044[22] << 44) +
      (src044[23] << 44) +
      (src044[24] << 44) +
      (src044[25] << 44) +
      (src044[26] << 44) +
      (src044[27] << 44) +
      (src044[28] << 44) +
      (src044[29] << 44) +
      (src044[30] << 44) +
      (src044[31] << 44) +
      (src044[32] << 44) +
      (src044[33] << 44) +
      (src044[34] << 44) +
      (src044[35] << 44) +
      (src044[36] << 44) +
      (src044[37] << 44) +
      (src044[38] << 44) +
      (src044[39] << 44) +
      (src044[40] << 44) +
      (src044[41] << 44) +
      (src044[42] << 44) +
      (src044[43] << 44) +
      (src044[44] << 44) +
      (src044[45] << 44) +
      (src044[46] << 44) +
      (src044[47] << 44) +
      (src044[48] << 44) +
      (src044[49] << 44) +
      (src044[50] << 44) +
      (src044[51] << 44) +
      (src044[52] << 44) +
      (src044[53] << 44) +
      (src044[54] << 44) +
      (src044[55] << 44) +
      (src044[56] << 44) +
      (src044[57] << 44) +
      (src044[58] << 44) +
      (src044[59] << 44) +
      (src044[60] << 44) +
      (src044[61] << 44) +
      (src044[62] << 44) +
      (src044[63] << 44) +
      (src044[64] << 44) +
      (src044[65] << 44) +
      (src044[66] << 44) +
      (src044[67] << 44) +
      (src044[68] << 44) +
      (src044[69] << 44) +
      (src044[70] << 44) +
      (src044[71] << 44) +
      (src044[72] << 44) +
      (src044[73] << 44) +
      (src044[74] << 44) +
      (src044[75] << 44) +
      (src044[76] << 44) +
      (src044[77] << 44) +
      (src044[78] << 44) +
      (src044[79] << 44) +
      (src044[80] << 44) +
      (src044[81] << 44) +
      (src044[82] << 44) +
      (src044[83] << 44) +
      (src044[84] << 44) +
      (src044[85] << 44) +
      (src044[86] << 44) +
      (src044[87] << 44) +
      (src044[88] << 44) +
      (src044[89] << 44) +
      (src044[90] << 44) +
      (src044[91] << 44) +
      (src044[92] << 44) +
      (src044[93] << 44) +
      (src044[94] << 44) +
      (src044[95] << 44) +
      (src044[96] << 44) +
      (src044[97] << 44) +
      (src044[98] << 44) +
      (src044[99] << 44) +
      (src044[100] << 44) +
      (src044[101] << 44) +
      (src044[102] << 44) +
      (src044[103] << 44) +
      (src044[104] << 44) +
      (src044[105] << 44) +
      (src044[106] << 44) +
      (src044[107] << 44) +
      (src044[108] << 44) +
      (src044[109] << 44) +
      (src044[110] << 44) +
      (src044[111] << 44) +
      (src044[112] << 44) +
      (src044[113] << 44) +
      (src044[114] << 44) +
      (src044[115] << 44) +
      (src044[116] << 44) +
      (src044[117] << 44) +
      (src044[118] << 44) +
      (src044[119] << 44) +
      (src044[120] << 44) +
      (src044[121] << 44) +
      (src044[122] << 44) +
      (src044[123] << 44) +
      (src044[124] << 44) +
      (src044[125] << 44) +
      (src044[126] << 44) +
      (src044[127] << 44) +
      (src045[0] << 45) +
      (src045[1] << 45) +
      (src045[2] << 45) +
      (src045[3] << 45) +
      (src045[4] << 45) +
      (src045[5] << 45) +
      (src045[6] << 45) +
      (src045[7] << 45) +
      (src045[8] << 45) +
      (src045[9] << 45) +
      (src045[10] << 45) +
      (src045[11] << 45) +
      (src045[12] << 45) +
      (src045[13] << 45) +
      (src045[14] << 45) +
      (src045[15] << 45) +
      (src045[16] << 45) +
      (src045[17] << 45) +
      (src045[18] << 45) +
      (src045[19] << 45) +
      (src045[20] << 45) +
      (src045[21] << 45) +
      (src045[22] << 45) +
      (src045[23] << 45) +
      (src045[24] << 45) +
      (src045[25] << 45) +
      (src045[26] << 45) +
      (src045[27] << 45) +
      (src045[28] << 45) +
      (src045[29] << 45) +
      (src045[30] << 45) +
      (src045[31] << 45) +
      (src045[32] << 45) +
      (src045[33] << 45) +
      (src045[34] << 45) +
      (src045[35] << 45) +
      (src045[36] << 45) +
      (src045[37] << 45) +
      (src045[38] << 45) +
      (src045[39] << 45) +
      (src045[40] << 45) +
      (src045[41] << 45) +
      (src045[42] << 45) +
      (src045[43] << 45) +
      (src045[44] << 45) +
      (src045[45] << 45) +
      (src045[46] << 45) +
      (src045[47] << 45) +
      (src045[48] << 45) +
      (src045[49] << 45) +
      (src045[50] << 45) +
      (src045[51] << 45) +
      (src045[52] << 45) +
      (src045[53] << 45) +
      (src045[54] << 45) +
      (src045[55] << 45) +
      (src045[56] << 45) +
      (src045[57] << 45) +
      (src045[58] << 45) +
      (src045[59] << 45) +
      (src045[60] << 45) +
      (src045[61] << 45) +
      (src045[62] << 45) +
      (src045[63] << 45) +
      (src045[64] << 45) +
      (src045[65] << 45) +
      (src045[66] << 45) +
      (src045[67] << 45) +
      (src045[68] << 45) +
      (src045[69] << 45) +
      (src045[70] << 45) +
      (src045[71] << 45) +
      (src045[72] << 45) +
      (src045[73] << 45) +
      (src045[74] << 45) +
      (src045[75] << 45) +
      (src045[76] << 45) +
      (src045[77] << 45) +
      (src045[78] << 45) +
      (src045[79] << 45) +
      (src045[80] << 45) +
      (src045[81] << 45) +
      (src045[82] << 45) +
      (src045[83] << 45) +
      (src045[84] << 45) +
      (src045[85] << 45) +
      (src045[86] << 45) +
      (src045[87] << 45) +
      (src045[88] << 45) +
      (src045[89] << 45) +
      (src045[90] << 45) +
      (src045[91] << 45) +
      (src045[92] << 45) +
      (src045[93] << 45) +
      (src045[94] << 45) +
      (src045[95] << 45) +
      (src045[96] << 45) +
      (src045[97] << 45) +
      (src045[98] << 45) +
      (src045[99] << 45) +
      (src045[100] << 45) +
      (src045[101] << 45) +
      (src045[102] << 45) +
      (src045[103] << 45) +
      (src045[104] << 45) +
      (src045[105] << 45) +
      (src045[106] << 45) +
      (src045[107] << 45) +
      (src045[108] << 45) +
      (src045[109] << 45) +
      (src045[110] << 45) +
      (src045[111] << 45) +
      (src045[112] << 45) +
      (src045[113] << 45) +
      (src045[114] << 45) +
      (src045[115] << 45) +
      (src045[116] << 45) +
      (src045[117] << 45) +
      (src045[118] << 45) +
      (src045[119] << 45) +
      (src045[120] << 45) +
      (src045[121] << 45) +
      (src045[122] << 45) +
      (src045[123] << 45) +
      (src045[124] << 45) +
      (src045[125] << 45) +
      (src045[126] << 45) +
      (src045[127] << 45) +
      (src046[0] << 46) +
      (src046[1] << 46) +
      (src046[2] << 46) +
      (src046[3] << 46) +
      (src046[4] << 46) +
      (src046[5] << 46) +
      (src046[6] << 46) +
      (src046[7] << 46) +
      (src046[8] << 46) +
      (src046[9] << 46) +
      (src046[10] << 46) +
      (src046[11] << 46) +
      (src046[12] << 46) +
      (src046[13] << 46) +
      (src046[14] << 46) +
      (src046[15] << 46) +
      (src046[16] << 46) +
      (src046[17] << 46) +
      (src046[18] << 46) +
      (src046[19] << 46) +
      (src046[20] << 46) +
      (src046[21] << 46) +
      (src046[22] << 46) +
      (src046[23] << 46) +
      (src046[24] << 46) +
      (src046[25] << 46) +
      (src046[26] << 46) +
      (src046[27] << 46) +
      (src046[28] << 46) +
      (src046[29] << 46) +
      (src046[30] << 46) +
      (src046[31] << 46) +
      (src046[32] << 46) +
      (src046[33] << 46) +
      (src046[34] << 46) +
      (src046[35] << 46) +
      (src046[36] << 46) +
      (src046[37] << 46) +
      (src046[38] << 46) +
      (src046[39] << 46) +
      (src046[40] << 46) +
      (src046[41] << 46) +
      (src046[42] << 46) +
      (src046[43] << 46) +
      (src046[44] << 46) +
      (src046[45] << 46) +
      (src046[46] << 46) +
      (src046[47] << 46) +
      (src046[48] << 46) +
      (src046[49] << 46) +
      (src046[50] << 46) +
      (src046[51] << 46) +
      (src046[52] << 46) +
      (src046[53] << 46) +
      (src046[54] << 46) +
      (src046[55] << 46) +
      (src046[56] << 46) +
      (src046[57] << 46) +
      (src046[58] << 46) +
      (src046[59] << 46) +
      (src046[60] << 46) +
      (src046[61] << 46) +
      (src046[62] << 46) +
      (src046[63] << 46) +
      (src046[64] << 46) +
      (src046[65] << 46) +
      (src046[66] << 46) +
      (src046[67] << 46) +
      (src046[68] << 46) +
      (src046[69] << 46) +
      (src046[70] << 46) +
      (src046[71] << 46) +
      (src046[72] << 46) +
      (src046[73] << 46) +
      (src046[74] << 46) +
      (src046[75] << 46) +
      (src046[76] << 46) +
      (src046[77] << 46) +
      (src046[78] << 46) +
      (src046[79] << 46) +
      (src046[80] << 46) +
      (src046[81] << 46) +
      (src046[82] << 46) +
      (src046[83] << 46) +
      (src046[84] << 46) +
      (src046[85] << 46) +
      (src046[86] << 46) +
      (src046[87] << 46) +
      (src046[88] << 46) +
      (src046[89] << 46) +
      (src046[90] << 46) +
      (src046[91] << 46) +
      (src046[92] << 46) +
      (src046[93] << 46) +
      (src046[94] << 46) +
      (src046[95] << 46) +
      (src046[96] << 46) +
      (src046[97] << 46) +
      (src046[98] << 46) +
      (src046[99] << 46) +
      (src046[100] << 46) +
      (src046[101] << 46) +
      (src046[102] << 46) +
      (src046[103] << 46) +
      (src046[104] << 46) +
      (src046[105] << 46) +
      (src046[106] << 46) +
      (src046[107] << 46) +
      (src046[108] << 46) +
      (src046[109] << 46) +
      (src046[110] << 46) +
      (src046[111] << 46) +
      (src046[112] << 46) +
      (src046[113] << 46) +
      (src046[114] << 46) +
      (src046[115] << 46) +
      (src046[116] << 46) +
      (src046[117] << 46) +
      (src046[118] << 46) +
      (src046[119] << 46) +
      (src046[120] << 46) +
      (src046[121] << 46) +
      (src046[122] << 46) +
      (src046[123] << 46) +
      (src046[124] << 46) +
      (src046[125] << 46) +
      (src046[126] << 46) +
      (src046[127] << 46) +
      (src047[0] << 47) +
      (src047[1] << 47) +
      (src047[2] << 47) +
      (src047[3] << 47) +
      (src047[4] << 47) +
      (src047[5] << 47) +
      (src047[6] << 47) +
      (src047[7] << 47) +
      (src047[8] << 47) +
      (src047[9] << 47) +
      (src047[10] << 47) +
      (src047[11] << 47) +
      (src047[12] << 47) +
      (src047[13] << 47) +
      (src047[14] << 47) +
      (src047[15] << 47) +
      (src047[16] << 47) +
      (src047[17] << 47) +
      (src047[18] << 47) +
      (src047[19] << 47) +
      (src047[20] << 47) +
      (src047[21] << 47) +
      (src047[22] << 47) +
      (src047[23] << 47) +
      (src047[24] << 47) +
      (src047[25] << 47) +
      (src047[26] << 47) +
      (src047[27] << 47) +
      (src047[28] << 47) +
      (src047[29] << 47) +
      (src047[30] << 47) +
      (src047[31] << 47) +
      (src047[32] << 47) +
      (src047[33] << 47) +
      (src047[34] << 47) +
      (src047[35] << 47) +
      (src047[36] << 47) +
      (src047[37] << 47) +
      (src047[38] << 47) +
      (src047[39] << 47) +
      (src047[40] << 47) +
      (src047[41] << 47) +
      (src047[42] << 47) +
      (src047[43] << 47) +
      (src047[44] << 47) +
      (src047[45] << 47) +
      (src047[46] << 47) +
      (src047[47] << 47) +
      (src047[48] << 47) +
      (src047[49] << 47) +
      (src047[50] << 47) +
      (src047[51] << 47) +
      (src047[52] << 47) +
      (src047[53] << 47) +
      (src047[54] << 47) +
      (src047[55] << 47) +
      (src047[56] << 47) +
      (src047[57] << 47) +
      (src047[58] << 47) +
      (src047[59] << 47) +
      (src047[60] << 47) +
      (src047[61] << 47) +
      (src047[62] << 47) +
      (src047[63] << 47) +
      (src047[64] << 47) +
      (src047[65] << 47) +
      (src047[66] << 47) +
      (src047[67] << 47) +
      (src047[68] << 47) +
      (src047[69] << 47) +
      (src047[70] << 47) +
      (src047[71] << 47) +
      (src047[72] << 47) +
      (src047[73] << 47) +
      (src047[74] << 47) +
      (src047[75] << 47) +
      (src047[76] << 47) +
      (src047[77] << 47) +
      (src047[78] << 47) +
      (src047[79] << 47) +
      (src047[80] << 47) +
      (src047[81] << 47) +
      (src047[82] << 47) +
      (src047[83] << 47) +
      (src047[84] << 47) +
      (src047[85] << 47) +
      (src047[86] << 47) +
      (src047[87] << 47) +
      (src047[88] << 47) +
      (src047[89] << 47) +
      (src047[90] << 47) +
      (src047[91] << 47) +
      (src047[92] << 47) +
      (src047[93] << 47) +
      (src047[94] << 47) +
      (src047[95] << 47) +
      (src047[96] << 47) +
      (src047[97] << 47) +
      (src047[98] << 47) +
      (src047[99] << 47) +
      (src047[100] << 47) +
      (src047[101] << 47) +
      (src047[102] << 47) +
      (src047[103] << 47) +
      (src047[104] << 47) +
      (src047[105] << 47) +
      (src047[106] << 47) +
      (src047[107] << 47) +
      (src047[108] << 47) +
      (src047[109] << 47) +
      (src047[110] << 47) +
      (src047[111] << 47) +
      (src047[112] << 47) +
      (src047[113] << 47) +
      (src047[114] << 47) +
      (src047[115] << 47) +
      (src047[116] << 47) +
      (src047[117] << 47) +
      (src047[118] << 47) +
      (src047[119] << 47) +
      (src047[120] << 47) +
      (src047[121] << 47) +
      (src047[122] << 47) +
      (src047[123] << 47) +
      (src047[124] << 47) +
      (src047[125] << 47) +
      (src047[126] << 47) +
      (src047[127] << 47) +
      (src048[0] << 48) +
      (src048[1] << 48) +
      (src048[2] << 48) +
      (src048[3] << 48) +
      (src048[4] << 48) +
      (src048[5] << 48) +
      (src048[6] << 48) +
      (src048[7] << 48) +
      (src048[8] << 48) +
      (src048[9] << 48) +
      (src048[10] << 48) +
      (src048[11] << 48) +
      (src048[12] << 48) +
      (src048[13] << 48) +
      (src048[14] << 48) +
      (src048[15] << 48) +
      (src048[16] << 48) +
      (src048[17] << 48) +
      (src048[18] << 48) +
      (src048[19] << 48) +
      (src048[20] << 48) +
      (src048[21] << 48) +
      (src048[22] << 48) +
      (src048[23] << 48) +
      (src048[24] << 48) +
      (src048[25] << 48) +
      (src048[26] << 48) +
      (src048[27] << 48) +
      (src048[28] << 48) +
      (src048[29] << 48) +
      (src048[30] << 48) +
      (src048[31] << 48) +
      (src048[32] << 48) +
      (src048[33] << 48) +
      (src048[34] << 48) +
      (src048[35] << 48) +
      (src048[36] << 48) +
      (src048[37] << 48) +
      (src048[38] << 48) +
      (src048[39] << 48) +
      (src048[40] << 48) +
      (src048[41] << 48) +
      (src048[42] << 48) +
      (src048[43] << 48) +
      (src048[44] << 48) +
      (src048[45] << 48) +
      (src048[46] << 48) +
      (src048[47] << 48) +
      (src048[48] << 48) +
      (src048[49] << 48) +
      (src048[50] << 48) +
      (src048[51] << 48) +
      (src048[52] << 48) +
      (src048[53] << 48) +
      (src048[54] << 48) +
      (src048[55] << 48) +
      (src048[56] << 48) +
      (src048[57] << 48) +
      (src048[58] << 48) +
      (src048[59] << 48) +
      (src048[60] << 48) +
      (src048[61] << 48) +
      (src048[62] << 48) +
      (src048[63] << 48) +
      (src048[64] << 48) +
      (src048[65] << 48) +
      (src048[66] << 48) +
      (src048[67] << 48) +
      (src048[68] << 48) +
      (src048[69] << 48) +
      (src048[70] << 48) +
      (src048[71] << 48) +
      (src048[72] << 48) +
      (src048[73] << 48) +
      (src048[74] << 48) +
      (src048[75] << 48) +
      (src048[76] << 48) +
      (src048[77] << 48) +
      (src048[78] << 48) +
      (src048[79] << 48) +
      (src048[80] << 48) +
      (src048[81] << 48) +
      (src048[82] << 48) +
      (src048[83] << 48) +
      (src048[84] << 48) +
      (src048[85] << 48) +
      (src048[86] << 48) +
      (src048[87] << 48) +
      (src048[88] << 48) +
      (src048[89] << 48) +
      (src048[90] << 48) +
      (src048[91] << 48) +
      (src048[92] << 48) +
      (src048[93] << 48) +
      (src048[94] << 48) +
      (src048[95] << 48) +
      (src048[96] << 48) +
      (src048[97] << 48) +
      (src048[98] << 48) +
      (src048[99] << 48) +
      (src048[100] << 48) +
      (src048[101] << 48) +
      (src048[102] << 48) +
      (src048[103] << 48) +
      (src048[104] << 48) +
      (src048[105] << 48) +
      (src048[106] << 48) +
      (src048[107] << 48) +
      (src048[108] << 48) +
      (src048[109] << 48) +
      (src048[110] << 48) +
      (src048[111] << 48) +
      (src048[112] << 48) +
      (src048[113] << 48) +
      (src048[114] << 48) +
      (src048[115] << 48) +
      (src048[116] << 48) +
      (src048[117] << 48) +
      (src048[118] << 48) +
      (src048[119] << 48) +
      (src048[120] << 48) +
      (src048[121] << 48) +
      (src048[122] << 48) +
      (src048[123] << 48) +
      (src048[124] << 48) +
      (src048[125] << 48) +
      (src048[126] << 48) +
      (src048[127] << 48) +
      (src049[0] << 49) +
      (src049[1] << 49) +
      (src049[2] << 49) +
      (src049[3] << 49) +
      (src049[4] << 49) +
      (src049[5] << 49) +
      (src049[6] << 49) +
      (src049[7] << 49) +
      (src049[8] << 49) +
      (src049[9] << 49) +
      (src049[10] << 49) +
      (src049[11] << 49) +
      (src049[12] << 49) +
      (src049[13] << 49) +
      (src049[14] << 49) +
      (src049[15] << 49) +
      (src049[16] << 49) +
      (src049[17] << 49) +
      (src049[18] << 49) +
      (src049[19] << 49) +
      (src049[20] << 49) +
      (src049[21] << 49) +
      (src049[22] << 49) +
      (src049[23] << 49) +
      (src049[24] << 49) +
      (src049[25] << 49) +
      (src049[26] << 49) +
      (src049[27] << 49) +
      (src049[28] << 49) +
      (src049[29] << 49) +
      (src049[30] << 49) +
      (src049[31] << 49) +
      (src049[32] << 49) +
      (src049[33] << 49) +
      (src049[34] << 49) +
      (src049[35] << 49) +
      (src049[36] << 49) +
      (src049[37] << 49) +
      (src049[38] << 49) +
      (src049[39] << 49) +
      (src049[40] << 49) +
      (src049[41] << 49) +
      (src049[42] << 49) +
      (src049[43] << 49) +
      (src049[44] << 49) +
      (src049[45] << 49) +
      (src049[46] << 49) +
      (src049[47] << 49) +
      (src049[48] << 49) +
      (src049[49] << 49) +
      (src049[50] << 49) +
      (src049[51] << 49) +
      (src049[52] << 49) +
      (src049[53] << 49) +
      (src049[54] << 49) +
      (src049[55] << 49) +
      (src049[56] << 49) +
      (src049[57] << 49) +
      (src049[58] << 49) +
      (src049[59] << 49) +
      (src049[60] << 49) +
      (src049[61] << 49) +
      (src049[62] << 49) +
      (src049[63] << 49) +
      (src049[64] << 49) +
      (src049[65] << 49) +
      (src049[66] << 49) +
      (src049[67] << 49) +
      (src049[68] << 49) +
      (src049[69] << 49) +
      (src049[70] << 49) +
      (src049[71] << 49) +
      (src049[72] << 49) +
      (src049[73] << 49) +
      (src049[74] << 49) +
      (src049[75] << 49) +
      (src049[76] << 49) +
      (src049[77] << 49) +
      (src049[78] << 49) +
      (src049[79] << 49) +
      (src049[80] << 49) +
      (src049[81] << 49) +
      (src049[82] << 49) +
      (src049[83] << 49) +
      (src049[84] << 49) +
      (src049[85] << 49) +
      (src049[86] << 49) +
      (src049[87] << 49) +
      (src049[88] << 49) +
      (src049[89] << 49) +
      (src049[90] << 49) +
      (src049[91] << 49) +
      (src049[92] << 49) +
      (src049[93] << 49) +
      (src049[94] << 49) +
      (src049[95] << 49) +
      (src049[96] << 49) +
      (src049[97] << 49) +
      (src049[98] << 49) +
      (src049[99] << 49) +
      (src049[100] << 49) +
      (src049[101] << 49) +
      (src049[102] << 49) +
      (src049[103] << 49) +
      (src049[104] << 49) +
      (src049[105] << 49) +
      (src049[106] << 49) +
      (src049[107] << 49) +
      (src049[108] << 49) +
      (src049[109] << 49) +
      (src049[110] << 49) +
      (src049[111] << 49) +
      (src049[112] << 49) +
      (src049[113] << 49) +
      (src049[114] << 49) +
      (src049[115] << 49) +
      (src049[116] << 49) +
      (src049[117] << 49) +
      (src049[118] << 49) +
      (src049[119] << 49) +
      (src049[120] << 49) +
      (src049[121] << 49) +
      (src049[122] << 49) +
      (src049[123] << 49) +
      (src049[124] << 49) +
      (src049[125] << 49) +
      (src049[126] << 49) +
      (src049[127] << 49) +
      (src050[0] << 50) +
      (src050[1] << 50) +
      (src050[2] << 50) +
      (src050[3] << 50) +
      (src050[4] << 50) +
      (src050[5] << 50) +
      (src050[6] << 50) +
      (src050[7] << 50) +
      (src050[8] << 50) +
      (src050[9] << 50) +
      (src050[10] << 50) +
      (src050[11] << 50) +
      (src050[12] << 50) +
      (src050[13] << 50) +
      (src050[14] << 50) +
      (src050[15] << 50) +
      (src050[16] << 50) +
      (src050[17] << 50) +
      (src050[18] << 50) +
      (src050[19] << 50) +
      (src050[20] << 50) +
      (src050[21] << 50) +
      (src050[22] << 50) +
      (src050[23] << 50) +
      (src050[24] << 50) +
      (src050[25] << 50) +
      (src050[26] << 50) +
      (src050[27] << 50) +
      (src050[28] << 50) +
      (src050[29] << 50) +
      (src050[30] << 50) +
      (src050[31] << 50) +
      (src050[32] << 50) +
      (src050[33] << 50) +
      (src050[34] << 50) +
      (src050[35] << 50) +
      (src050[36] << 50) +
      (src050[37] << 50) +
      (src050[38] << 50) +
      (src050[39] << 50) +
      (src050[40] << 50) +
      (src050[41] << 50) +
      (src050[42] << 50) +
      (src050[43] << 50) +
      (src050[44] << 50) +
      (src050[45] << 50) +
      (src050[46] << 50) +
      (src050[47] << 50) +
      (src050[48] << 50) +
      (src050[49] << 50) +
      (src050[50] << 50) +
      (src050[51] << 50) +
      (src050[52] << 50) +
      (src050[53] << 50) +
      (src050[54] << 50) +
      (src050[55] << 50) +
      (src050[56] << 50) +
      (src050[57] << 50) +
      (src050[58] << 50) +
      (src050[59] << 50) +
      (src050[60] << 50) +
      (src050[61] << 50) +
      (src050[62] << 50) +
      (src050[63] << 50) +
      (src050[64] << 50) +
      (src050[65] << 50) +
      (src050[66] << 50) +
      (src050[67] << 50) +
      (src050[68] << 50) +
      (src050[69] << 50) +
      (src050[70] << 50) +
      (src050[71] << 50) +
      (src050[72] << 50) +
      (src050[73] << 50) +
      (src050[74] << 50) +
      (src050[75] << 50) +
      (src050[76] << 50) +
      (src050[77] << 50) +
      (src050[78] << 50) +
      (src050[79] << 50) +
      (src050[80] << 50) +
      (src050[81] << 50) +
      (src050[82] << 50) +
      (src050[83] << 50) +
      (src050[84] << 50) +
      (src050[85] << 50) +
      (src050[86] << 50) +
      (src050[87] << 50) +
      (src050[88] << 50) +
      (src050[89] << 50) +
      (src050[90] << 50) +
      (src050[91] << 50) +
      (src050[92] << 50) +
      (src050[93] << 50) +
      (src050[94] << 50) +
      (src050[95] << 50) +
      (src050[96] << 50) +
      (src050[97] << 50) +
      (src050[98] << 50) +
      (src050[99] << 50) +
      (src050[100] << 50) +
      (src050[101] << 50) +
      (src050[102] << 50) +
      (src050[103] << 50) +
      (src050[104] << 50) +
      (src050[105] << 50) +
      (src050[106] << 50) +
      (src050[107] << 50) +
      (src050[108] << 50) +
      (src050[109] << 50) +
      (src050[110] << 50) +
      (src050[111] << 50) +
      (src050[112] << 50) +
      (src050[113] << 50) +
      (src050[114] << 50) +
      (src050[115] << 50) +
      (src050[116] << 50) +
      (src050[117] << 50) +
      (src050[118] << 50) +
      (src050[119] << 50) +
      (src050[120] << 50) +
      (src050[121] << 50) +
      (src050[122] << 50) +
      (src050[123] << 50) +
      (src050[124] << 50) +
      (src050[125] << 50) +
      (src050[126] << 50) +
      (src050[127] << 50) +
      (src051[0] << 51) +
      (src051[1] << 51) +
      (src051[2] << 51) +
      (src051[3] << 51) +
      (src051[4] << 51) +
      (src051[5] << 51) +
      (src051[6] << 51) +
      (src051[7] << 51) +
      (src051[8] << 51) +
      (src051[9] << 51) +
      (src051[10] << 51) +
      (src051[11] << 51) +
      (src051[12] << 51) +
      (src051[13] << 51) +
      (src051[14] << 51) +
      (src051[15] << 51) +
      (src051[16] << 51) +
      (src051[17] << 51) +
      (src051[18] << 51) +
      (src051[19] << 51) +
      (src051[20] << 51) +
      (src051[21] << 51) +
      (src051[22] << 51) +
      (src051[23] << 51) +
      (src051[24] << 51) +
      (src051[25] << 51) +
      (src051[26] << 51) +
      (src051[27] << 51) +
      (src051[28] << 51) +
      (src051[29] << 51) +
      (src051[30] << 51) +
      (src051[31] << 51) +
      (src051[32] << 51) +
      (src051[33] << 51) +
      (src051[34] << 51) +
      (src051[35] << 51) +
      (src051[36] << 51) +
      (src051[37] << 51) +
      (src051[38] << 51) +
      (src051[39] << 51) +
      (src051[40] << 51) +
      (src051[41] << 51) +
      (src051[42] << 51) +
      (src051[43] << 51) +
      (src051[44] << 51) +
      (src051[45] << 51) +
      (src051[46] << 51) +
      (src051[47] << 51) +
      (src051[48] << 51) +
      (src051[49] << 51) +
      (src051[50] << 51) +
      (src051[51] << 51) +
      (src051[52] << 51) +
      (src051[53] << 51) +
      (src051[54] << 51) +
      (src051[55] << 51) +
      (src051[56] << 51) +
      (src051[57] << 51) +
      (src051[58] << 51) +
      (src051[59] << 51) +
      (src051[60] << 51) +
      (src051[61] << 51) +
      (src051[62] << 51) +
      (src051[63] << 51) +
      (src051[64] << 51) +
      (src051[65] << 51) +
      (src051[66] << 51) +
      (src051[67] << 51) +
      (src051[68] << 51) +
      (src051[69] << 51) +
      (src051[70] << 51) +
      (src051[71] << 51) +
      (src051[72] << 51) +
      (src051[73] << 51) +
      (src051[74] << 51) +
      (src051[75] << 51) +
      (src051[76] << 51) +
      (src051[77] << 51) +
      (src051[78] << 51) +
      (src051[79] << 51) +
      (src051[80] << 51) +
      (src051[81] << 51) +
      (src051[82] << 51) +
      (src051[83] << 51) +
      (src051[84] << 51) +
      (src051[85] << 51) +
      (src051[86] << 51) +
      (src051[87] << 51) +
      (src051[88] << 51) +
      (src051[89] << 51) +
      (src051[90] << 51) +
      (src051[91] << 51) +
      (src051[92] << 51) +
      (src051[93] << 51) +
      (src051[94] << 51) +
      (src051[95] << 51) +
      (src051[96] << 51) +
      (src051[97] << 51) +
      (src051[98] << 51) +
      (src051[99] << 51) +
      (src051[100] << 51) +
      (src051[101] << 51) +
      (src051[102] << 51) +
      (src051[103] << 51) +
      (src051[104] << 51) +
      (src051[105] << 51) +
      (src051[106] << 51) +
      (src051[107] << 51) +
      (src051[108] << 51) +
      (src051[109] << 51) +
      (src051[110] << 51) +
      (src051[111] << 51) +
      (src051[112] << 51) +
      (src051[113] << 51) +
      (src051[114] << 51) +
      (src051[115] << 51) +
      (src051[116] << 51) +
      (src051[117] << 51) +
      (src051[118] << 51) +
      (src051[119] << 51) +
      (src051[120] << 51) +
      (src051[121] << 51) +
      (src051[122] << 51) +
      (src051[123] << 51) +
      (src051[124] << 51) +
      (src051[125] << 51) +
      (src051[126] << 51) +
      (src051[127] << 51) +
      (src052[0] << 52) +
      (src052[1] << 52) +
      (src052[2] << 52) +
      (src052[3] << 52) +
      (src052[4] << 52) +
      (src052[5] << 52) +
      (src052[6] << 52) +
      (src052[7] << 52) +
      (src052[8] << 52) +
      (src052[9] << 52) +
      (src052[10] << 52) +
      (src052[11] << 52) +
      (src052[12] << 52) +
      (src052[13] << 52) +
      (src052[14] << 52) +
      (src052[15] << 52) +
      (src052[16] << 52) +
      (src052[17] << 52) +
      (src052[18] << 52) +
      (src052[19] << 52) +
      (src052[20] << 52) +
      (src052[21] << 52) +
      (src052[22] << 52) +
      (src052[23] << 52) +
      (src052[24] << 52) +
      (src052[25] << 52) +
      (src052[26] << 52) +
      (src052[27] << 52) +
      (src052[28] << 52) +
      (src052[29] << 52) +
      (src052[30] << 52) +
      (src052[31] << 52) +
      (src052[32] << 52) +
      (src052[33] << 52) +
      (src052[34] << 52) +
      (src052[35] << 52) +
      (src052[36] << 52) +
      (src052[37] << 52) +
      (src052[38] << 52) +
      (src052[39] << 52) +
      (src052[40] << 52) +
      (src052[41] << 52) +
      (src052[42] << 52) +
      (src052[43] << 52) +
      (src052[44] << 52) +
      (src052[45] << 52) +
      (src052[46] << 52) +
      (src052[47] << 52) +
      (src052[48] << 52) +
      (src052[49] << 52) +
      (src052[50] << 52) +
      (src052[51] << 52) +
      (src052[52] << 52) +
      (src052[53] << 52) +
      (src052[54] << 52) +
      (src052[55] << 52) +
      (src052[56] << 52) +
      (src052[57] << 52) +
      (src052[58] << 52) +
      (src052[59] << 52) +
      (src052[60] << 52) +
      (src052[61] << 52) +
      (src052[62] << 52) +
      (src052[63] << 52) +
      (src052[64] << 52) +
      (src052[65] << 52) +
      (src052[66] << 52) +
      (src052[67] << 52) +
      (src052[68] << 52) +
      (src052[69] << 52) +
      (src052[70] << 52) +
      (src052[71] << 52) +
      (src052[72] << 52) +
      (src052[73] << 52) +
      (src052[74] << 52) +
      (src052[75] << 52) +
      (src052[76] << 52) +
      (src052[77] << 52) +
      (src052[78] << 52) +
      (src052[79] << 52) +
      (src052[80] << 52) +
      (src052[81] << 52) +
      (src052[82] << 52) +
      (src052[83] << 52) +
      (src052[84] << 52) +
      (src052[85] << 52) +
      (src052[86] << 52) +
      (src052[87] << 52) +
      (src052[88] << 52) +
      (src052[89] << 52) +
      (src052[90] << 52) +
      (src052[91] << 52) +
      (src052[92] << 52) +
      (src052[93] << 52) +
      (src052[94] << 52) +
      (src052[95] << 52) +
      (src052[96] << 52) +
      (src052[97] << 52) +
      (src052[98] << 52) +
      (src052[99] << 52) +
      (src052[100] << 52) +
      (src052[101] << 52) +
      (src052[102] << 52) +
      (src052[103] << 52) +
      (src052[104] << 52) +
      (src052[105] << 52) +
      (src052[106] << 52) +
      (src052[107] << 52) +
      (src052[108] << 52) +
      (src052[109] << 52) +
      (src052[110] << 52) +
      (src052[111] << 52) +
      (src052[112] << 52) +
      (src052[113] << 52) +
      (src052[114] << 52) +
      (src052[115] << 52) +
      (src052[116] << 52) +
      (src052[117] << 52) +
      (src052[118] << 52) +
      (src052[119] << 52) +
      (src052[120] << 52) +
      (src052[121] << 52) +
      (src052[122] << 52) +
      (src052[123] << 52) +
      (src052[124] << 52) +
      (src052[125] << 52) +
      (src052[126] << 52) +
      (src052[127] << 52) +
      (src053[0] << 53) +
      (src053[1] << 53) +
      (src053[2] << 53) +
      (src053[3] << 53) +
      (src053[4] << 53) +
      (src053[5] << 53) +
      (src053[6] << 53) +
      (src053[7] << 53) +
      (src053[8] << 53) +
      (src053[9] << 53) +
      (src053[10] << 53) +
      (src053[11] << 53) +
      (src053[12] << 53) +
      (src053[13] << 53) +
      (src053[14] << 53) +
      (src053[15] << 53) +
      (src053[16] << 53) +
      (src053[17] << 53) +
      (src053[18] << 53) +
      (src053[19] << 53) +
      (src053[20] << 53) +
      (src053[21] << 53) +
      (src053[22] << 53) +
      (src053[23] << 53) +
      (src053[24] << 53) +
      (src053[25] << 53) +
      (src053[26] << 53) +
      (src053[27] << 53) +
      (src053[28] << 53) +
      (src053[29] << 53) +
      (src053[30] << 53) +
      (src053[31] << 53) +
      (src053[32] << 53) +
      (src053[33] << 53) +
      (src053[34] << 53) +
      (src053[35] << 53) +
      (src053[36] << 53) +
      (src053[37] << 53) +
      (src053[38] << 53) +
      (src053[39] << 53) +
      (src053[40] << 53) +
      (src053[41] << 53) +
      (src053[42] << 53) +
      (src053[43] << 53) +
      (src053[44] << 53) +
      (src053[45] << 53) +
      (src053[46] << 53) +
      (src053[47] << 53) +
      (src053[48] << 53) +
      (src053[49] << 53) +
      (src053[50] << 53) +
      (src053[51] << 53) +
      (src053[52] << 53) +
      (src053[53] << 53) +
      (src053[54] << 53) +
      (src053[55] << 53) +
      (src053[56] << 53) +
      (src053[57] << 53) +
      (src053[58] << 53) +
      (src053[59] << 53) +
      (src053[60] << 53) +
      (src053[61] << 53) +
      (src053[62] << 53) +
      (src053[63] << 53) +
      (src053[64] << 53) +
      (src053[65] << 53) +
      (src053[66] << 53) +
      (src053[67] << 53) +
      (src053[68] << 53) +
      (src053[69] << 53) +
      (src053[70] << 53) +
      (src053[71] << 53) +
      (src053[72] << 53) +
      (src053[73] << 53) +
      (src053[74] << 53) +
      (src053[75] << 53) +
      (src053[76] << 53) +
      (src053[77] << 53) +
      (src053[78] << 53) +
      (src053[79] << 53) +
      (src053[80] << 53) +
      (src053[81] << 53) +
      (src053[82] << 53) +
      (src053[83] << 53) +
      (src053[84] << 53) +
      (src053[85] << 53) +
      (src053[86] << 53) +
      (src053[87] << 53) +
      (src053[88] << 53) +
      (src053[89] << 53) +
      (src053[90] << 53) +
      (src053[91] << 53) +
      (src053[92] << 53) +
      (src053[93] << 53) +
      (src053[94] << 53) +
      (src053[95] << 53) +
      (src053[96] << 53) +
      (src053[97] << 53) +
      (src053[98] << 53) +
      (src053[99] << 53) +
      (src053[100] << 53) +
      (src053[101] << 53) +
      (src053[102] << 53) +
      (src053[103] << 53) +
      (src053[104] << 53) +
      (src053[105] << 53) +
      (src053[106] << 53) +
      (src053[107] << 53) +
      (src053[108] << 53) +
      (src053[109] << 53) +
      (src053[110] << 53) +
      (src053[111] << 53) +
      (src053[112] << 53) +
      (src053[113] << 53) +
      (src053[114] << 53) +
      (src053[115] << 53) +
      (src053[116] << 53) +
      (src053[117] << 53) +
      (src053[118] << 53) +
      (src053[119] << 53) +
      (src053[120] << 53) +
      (src053[121] << 53) +
      (src053[122] << 53) +
      (src053[123] << 53) +
      (src053[124] << 53) +
      (src053[125] << 53) +
      (src053[126] << 53) +
      (src053[127] << 53) +
      (src054[0] << 54) +
      (src054[1] << 54) +
      (src054[2] << 54) +
      (src054[3] << 54) +
      (src054[4] << 54) +
      (src054[5] << 54) +
      (src054[6] << 54) +
      (src054[7] << 54) +
      (src054[8] << 54) +
      (src054[9] << 54) +
      (src054[10] << 54) +
      (src054[11] << 54) +
      (src054[12] << 54) +
      (src054[13] << 54) +
      (src054[14] << 54) +
      (src054[15] << 54) +
      (src054[16] << 54) +
      (src054[17] << 54) +
      (src054[18] << 54) +
      (src054[19] << 54) +
      (src054[20] << 54) +
      (src054[21] << 54) +
      (src054[22] << 54) +
      (src054[23] << 54) +
      (src054[24] << 54) +
      (src054[25] << 54) +
      (src054[26] << 54) +
      (src054[27] << 54) +
      (src054[28] << 54) +
      (src054[29] << 54) +
      (src054[30] << 54) +
      (src054[31] << 54) +
      (src054[32] << 54) +
      (src054[33] << 54) +
      (src054[34] << 54) +
      (src054[35] << 54) +
      (src054[36] << 54) +
      (src054[37] << 54) +
      (src054[38] << 54) +
      (src054[39] << 54) +
      (src054[40] << 54) +
      (src054[41] << 54) +
      (src054[42] << 54) +
      (src054[43] << 54) +
      (src054[44] << 54) +
      (src054[45] << 54) +
      (src054[46] << 54) +
      (src054[47] << 54) +
      (src054[48] << 54) +
      (src054[49] << 54) +
      (src054[50] << 54) +
      (src054[51] << 54) +
      (src054[52] << 54) +
      (src054[53] << 54) +
      (src054[54] << 54) +
      (src054[55] << 54) +
      (src054[56] << 54) +
      (src054[57] << 54) +
      (src054[58] << 54) +
      (src054[59] << 54) +
      (src054[60] << 54) +
      (src054[61] << 54) +
      (src054[62] << 54) +
      (src054[63] << 54) +
      (src054[64] << 54) +
      (src054[65] << 54) +
      (src054[66] << 54) +
      (src054[67] << 54) +
      (src054[68] << 54) +
      (src054[69] << 54) +
      (src054[70] << 54) +
      (src054[71] << 54) +
      (src054[72] << 54) +
      (src054[73] << 54) +
      (src054[74] << 54) +
      (src054[75] << 54) +
      (src054[76] << 54) +
      (src054[77] << 54) +
      (src054[78] << 54) +
      (src054[79] << 54) +
      (src054[80] << 54) +
      (src054[81] << 54) +
      (src054[82] << 54) +
      (src054[83] << 54) +
      (src054[84] << 54) +
      (src054[85] << 54) +
      (src054[86] << 54) +
      (src054[87] << 54) +
      (src054[88] << 54) +
      (src054[89] << 54) +
      (src054[90] << 54) +
      (src054[91] << 54) +
      (src054[92] << 54) +
      (src054[93] << 54) +
      (src054[94] << 54) +
      (src054[95] << 54) +
      (src054[96] << 54) +
      (src054[97] << 54) +
      (src054[98] << 54) +
      (src054[99] << 54) +
      (src054[100] << 54) +
      (src054[101] << 54) +
      (src054[102] << 54) +
      (src054[103] << 54) +
      (src054[104] << 54) +
      (src054[105] << 54) +
      (src054[106] << 54) +
      (src054[107] << 54) +
      (src054[108] << 54) +
      (src054[109] << 54) +
      (src054[110] << 54) +
      (src054[111] << 54) +
      (src054[112] << 54) +
      (src054[113] << 54) +
      (src054[114] << 54) +
      (src054[115] << 54) +
      (src054[116] << 54) +
      (src054[117] << 54) +
      (src054[118] << 54) +
      (src054[119] << 54) +
      (src054[120] << 54) +
      (src054[121] << 54) +
      (src054[122] << 54) +
      (src054[123] << 54) +
      (src054[124] << 54) +
      (src054[125] << 54) +
      (src054[126] << 54) +
      (src054[127] << 54) +
      (src055[0] << 55) +
      (src055[1] << 55) +
      (src055[2] << 55) +
      (src055[3] << 55) +
      (src055[4] << 55) +
      (src055[5] << 55) +
      (src055[6] << 55) +
      (src055[7] << 55) +
      (src055[8] << 55) +
      (src055[9] << 55) +
      (src055[10] << 55) +
      (src055[11] << 55) +
      (src055[12] << 55) +
      (src055[13] << 55) +
      (src055[14] << 55) +
      (src055[15] << 55) +
      (src055[16] << 55) +
      (src055[17] << 55) +
      (src055[18] << 55) +
      (src055[19] << 55) +
      (src055[20] << 55) +
      (src055[21] << 55) +
      (src055[22] << 55) +
      (src055[23] << 55) +
      (src055[24] << 55) +
      (src055[25] << 55) +
      (src055[26] << 55) +
      (src055[27] << 55) +
      (src055[28] << 55) +
      (src055[29] << 55) +
      (src055[30] << 55) +
      (src055[31] << 55) +
      (src055[32] << 55) +
      (src055[33] << 55) +
      (src055[34] << 55) +
      (src055[35] << 55) +
      (src055[36] << 55) +
      (src055[37] << 55) +
      (src055[38] << 55) +
      (src055[39] << 55) +
      (src055[40] << 55) +
      (src055[41] << 55) +
      (src055[42] << 55) +
      (src055[43] << 55) +
      (src055[44] << 55) +
      (src055[45] << 55) +
      (src055[46] << 55) +
      (src055[47] << 55) +
      (src055[48] << 55) +
      (src055[49] << 55) +
      (src055[50] << 55) +
      (src055[51] << 55) +
      (src055[52] << 55) +
      (src055[53] << 55) +
      (src055[54] << 55) +
      (src055[55] << 55) +
      (src055[56] << 55) +
      (src055[57] << 55) +
      (src055[58] << 55) +
      (src055[59] << 55) +
      (src055[60] << 55) +
      (src055[61] << 55) +
      (src055[62] << 55) +
      (src055[63] << 55) +
      (src055[64] << 55) +
      (src055[65] << 55) +
      (src055[66] << 55) +
      (src055[67] << 55) +
      (src055[68] << 55) +
      (src055[69] << 55) +
      (src055[70] << 55) +
      (src055[71] << 55) +
      (src055[72] << 55) +
      (src055[73] << 55) +
      (src055[74] << 55) +
      (src055[75] << 55) +
      (src055[76] << 55) +
      (src055[77] << 55) +
      (src055[78] << 55) +
      (src055[79] << 55) +
      (src055[80] << 55) +
      (src055[81] << 55) +
      (src055[82] << 55) +
      (src055[83] << 55) +
      (src055[84] << 55) +
      (src055[85] << 55) +
      (src055[86] << 55) +
      (src055[87] << 55) +
      (src055[88] << 55) +
      (src055[89] << 55) +
      (src055[90] << 55) +
      (src055[91] << 55) +
      (src055[92] << 55) +
      (src055[93] << 55) +
      (src055[94] << 55) +
      (src055[95] << 55) +
      (src055[96] << 55) +
      (src055[97] << 55) +
      (src055[98] << 55) +
      (src055[99] << 55) +
      (src055[100] << 55) +
      (src055[101] << 55) +
      (src055[102] << 55) +
      (src055[103] << 55) +
      (src055[104] << 55) +
      (src055[105] << 55) +
      (src055[106] << 55) +
      (src055[107] << 55) +
      (src055[108] << 55) +
      (src055[109] << 55) +
      (src055[110] << 55) +
      (src055[111] << 55) +
      (src055[112] << 55) +
      (src055[113] << 55) +
      (src055[114] << 55) +
      (src055[115] << 55) +
      (src055[116] << 55) +
      (src055[117] << 55) +
      (src055[118] << 55) +
      (src055[119] << 55) +
      (src055[120] << 55) +
      (src055[121] << 55) +
      (src055[122] << 55) +
      (src055[123] << 55) +
      (src055[124] << 55) +
      (src055[125] << 55) +
      (src055[126] << 55) +
      (src055[127] << 55) +
      (src056[0] << 56) +
      (src056[1] << 56) +
      (src056[2] << 56) +
      (src056[3] << 56) +
      (src056[4] << 56) +
      (src056[5] << 56) +
      (src056[6] << 56) +
      (src056[7] << 56) +
      (src056[8] << 56) +
      (src056[9] << 56) +
      (src056[10] << 56) +
      (src056[11] << 56) +
      (src056[12] << 56) +
      (src056[13] << 56) +
      (src056[14] << 56) +
      (src056[15] << 56) +
      (src056[16] << 56) +
      (src056[17] << 56) +
      (src056[18] << 56) +
      (src056[19] << 56) +
      (src056[20] << 56) +
      (src056[21] << 56) +
      (src056[22] << 56) +
      (src056[23] << 56) +
      (src056[24] << 56) +
      (src056[25] << 56) +
      (src056[26] << 56) +
      (src056[27] << 56) +
      (src056[28] << 56) +
      (src056[29] << 56) +
      (src056[30] << 56) +
      (src056[31] << 56) +
      (src056[32] << 56) +
      (src056[33] << 56) +
      (src056[34] << 56) +
      (src056[35] << 56) +
      (src056[36] << 56) +
      (src056[37] << 56) +
      (src056[38] << 56) +
      (src056[39] << 56) +
      (src056[40] << 56) +
      (src056[41] << 56) +
      (src056[42] << 56) +
      (src056[43] << 56) +
      (src056[44] << 56) +
      (src056[45] << 56) +
      (src056[46] << 56) +
      (src056[47] << 56) +
      (src056[48] << 56) +
      (src056[49] << 56) +
      (src056[50] << 56) +
      (src056[51] << 56) +
      (src056[52] << 56) +
      (src056[53] << 56) +
      (src056[54] << 56) +
      (src056[55] << 56) +
      (src056[56] << 56) +
      (src056[57] << 56) +
      (src056[58] << 56) +
      (src056[59] << 56) +
      (src056[60] << 56) +
      (src056[61] << 56) +
      (src056[62] << 56) +
      (src056[63] << 56) +
      (src056[64] << 56) +
      (src056[65] << 56) +
      (src056[66] << 56) +
      (src056[67] << 56) +
      (src056[68] << 56) +
      (src056[69] << 56) +
      (src056[70] << 56) +
      (src056[71] << 56) +
      (src056[72] << 56) +
      (src056[73] << 56) +
      (src056[74] << 56) +
      (src056[75] << 56) +
      (src056[76] << 56) +
      (src056[77] << 56) +
      (src056[78] << 56) +
      (src056[79] << 56) +
      (src056[80] << 56) +
      (src056[81] << 56) +
      (src056[82] << 56) +
      (src056[83] << 56) +
      (src056[84] << 56) +
      (src056[85] << 56) +
      (src056[86] << 56) +
      (src056[87] << 56) +
      (src056[88] << 56) +
      (src056[89] << 56) +
      (src056[90] << 56) +
      (src056[91] << 56) +
      (src056[92] << 56) +
      (src056[93] << 56) +
      (src056[94] << 56) +
      (src056[95] << 56) +
      (src056[96] << 56) +
      (src056[97] << 56) +
      (src056[98] << 56) +
      (src056[99] << 56) +
      (src056[100] << 56) +
      (src056[101] << 56) +
      (src056[102] << 56) +
      (src056[103] << 56) +
      (src056[104] << 56) +
      (src056[105] << 56) +
      (src056[106] << 56) +
      (src056[107] << 56) +
      (src056[108] << 56) +
      (src056[109] << 56) +
      (src056[110] << 56) +
      (src056[111] << 56) +
      (src056[112] << 56) +
      (src056[113] << 56) +
      (src056[114] << 56) +
      (src056[115] << 56) +
      (src056[116] << 56) +
      (src056[117] << 56) +
      (src056[118] << 56) +
      (src056[119] << 56) +
      (src056[120] << 56) +
      (src056[121] << 56) +
      (src056[122] << 56) +
      (src056[123] << 56) +
      (src056[124] << 56) +
      (src056[125] << 56) +
      (src056[126] << 56) +
      (src056[127] << 56) +
      (src057[0] << 57) +
      (src057[1] << 57) +
      (src057[2] << 57) +
      (src057[3] << 57) +
      (src057[4] << 57) +
      (src057[5] << 57) +
      (src057[6] << 57) +
      (src057[7] << 57) +
      (src057[8] << 57) +
      (src057[9] << 57) +
      (src057[10] << 57) +
      (src057[11] << 57) +
      (src057[12] << 57) +
      (src057[13] << 57) +
      (src057[14] << 57) +
      (src057[15] << 57) +
      (src057[16] << 57) +
      (src057[17] << 57) +
      (src057[18] << 57) +
      (src057[19] << 57) +
      (src057[20] << 57) +
      (src057[21] << 57) +
      (src057[22] << 57) +
      (src057[23] << 57) +
      (src057[24] << 57) +
      (src057[25] << 57) +
      (src057[26] << 57) +
      (src057[27] << 57) +
      (src057[28] << 57) +
      (src057[29] << 57) +
      (src057[30] << 57) +
      (src057[31] << 57) +
      (src057[32] << 57) +
      (src057[33] << 57) +
      (src057[34] << 57) +
      (src057[35] << 57) +
      (src057[36] << 57) +
      (src057[37] << 57) +
      (src057[38] << 57) +
      (src057[39] << 57) +
      (src057[40] << 57) +
      (src057[41] << 57) +
      (src057[42] << 57) +
      (src057[43] << 57) +
      (src057[44] << 57) +
      (src057[45] << 57) +
      (src057[46] << 57) +
      (src057[47] << 57) +
      (src057[48] << 57) +
      (src057[49] << 57) +
      (src057[50] << 57) +
      (src057[51] << 57) +
      (src057[52] << 57) +
      (src057[53] << 57) +
      (src057[54] << 57) +
      (src057[55] << 57) +
      (src057[56] << 57) +
      (src057[57] << 57) +
      (src057[58] << 57) +
      (src057[59] << 57) +
      (src057[60] << 57) +
      (src057[61] << 57) +
      (src057[62] << 57) +
      (src057[63] << 57) +
      (src057[64] << 57) +
      (src057[65] << 57) +
      (src057[66] << 57) +
      (src057[67] << 57) +
      (src057[68] << 57) +
      (src057[69] << 57) +
      (src057[70] << 57) +
      (src057[71] << 57) +
      (src057[72] << 57) +
      (src057[73] << 57) +
      (src057[74] << 57) +
      (src057[75] << 57) +
      (src057[76] << 57) +
      (src057[77] << 57) +
      (src057[78] << 57) +
      (src057[79] << 57) +
      (src057[80] << 57) +
      (src057[81] << 57) +
      (src057[82] << 57) +
      (src057[83] << 57) +
      (src057[84] << 57) +
      (src057[85] << 57) +
      (src057[86] << 57) +
      (src057[87] << 57) +
      (src057[88] << 57) +
      (src057[89] << 57) +
      (src057[90] << 57) +
      (src057[91] << 57) +
      (src057[92] << 57) +
      (src057[93] << 57) +
      (src057[94] << 57) +
      (src057[95] << 57) +
      (src057[96] << 57) +
      (src057[97] << 57) +
      (src057[98] << 57) +
      (src057[99] << 57) +
      (src057[100] << 57) +
      (src057[101] << 57) +
      (src057[102] << 57) +
      (src057[103] << 57) +
      (src057[104] << 57) +
      (src057[105] << 57) +
      (src057[106] << 57) +
      (src057[107] << 57) +
      (src057[108] << 57) +
      (src057[109] << 57) +
      (src057[110] << 57) +
      (src057[111] << 57) +
      (src057[112] << 57) +
      (src057[113] << 57) +
      (src057[114] << 57) +
      (src057[115] << 57) +
      (src057[116] << 57) +
      (src057[117] << 57) +
      (src057[118] << 57) +
      (src057[119] << 57) +
      (src057[120] << 57) +
      (src057[121] << 57) +
      (src057[122] << 57) +
      (src057[123] << 57) +
      (src057[124] << 57) +
      (src057[125] << 57) +
      (src057[126] << 57) +
      (src057[127] << 57) +
      (src058[0] << 58) +
      (src058[1] << 58) +
      (src058[2] << 58) +
      (src058[3] << 58) +
      (src058[4] << 58) +
      (src058[5] << 58) +
      (src058[6] << 58) +
      (src058[7] << 58) +
      (src058[8] << 58) +
      (src058[9] << 58) +
      (src058[10] << 58) +
      (src058[11] << 58) +
      (src058[12] << 58) +
      (src058[13] << 58) +
      (src058[14] << 58) +
      (src058[15] << 58) +
      (src058[16] << 58) +
      (src058[17] << 58) +
      (src058[18] << 58) +
      (src058[19] << 58) +
      (src058[20] << 58) +
      (src058[21] << 58) +
      (src058[22] << 58) +
      (src058[23] << 58) +
      (src058[24] << 58) +
      (src058[25] << 58) +
      (src058[26] << 58) +
      (src058[27] << 58) +
      (src058[28] << 58) +
      (src058[29] << 58) +
      (src058[30] << 58) +
      (src058[31] << 58) +
      (src058[32] << 58) +
      (src058[33] << 58) +
      (src058[34] << 58) +
      (src058[35] << 58) +
      (src058[36] << 58) +
      (src058[37] << 58) +
      (src058[38] << 58) +
      (src058[39] << 58) +
      (src058[40] << 58) +
      (src058[41] << 58) +
      (src058[42] << 58) +
      (src058[43] << 58) +
      (src058[44] << 58) +
      (src058[45] << 58) +
      (src058[46] << 58) +
      (src058[47] << 58) +
      (src058[48] << 58) +
      (src058[49] << 58) +
      (src058[50] << 58) +
      (src058[51] << 58) +
      (src058[52] << 58) +
      (src058[53] << 58) +
      (src058[54] << 58) +
      (src058[55] << 58) +
      (src058[56] << 58) +
      (src058[57] << 58) +
      (src058[58] << 58) +
      (src058[59] << 58) +
      (src058[60] << 58) +
      (src058[61] << 58) +
      (src058[62] << 58) +
      (src058[63] << 58) +
      (src058[64] << 58) +
      (src058[65] << 58) +
      (src058[66] << 58) +
      (src058[67] << 58) +
      (src058[68] << 58) +
      (src058[69] << 58) +
      (src058[70] << 58) +
      (src058[71] << 58) +
      (src058[72] << 58) +
      (src058[73] << 58) +
      (src058[74] << 58) +
      (src058[75] << 58) +
      (src058[76] << 58) +
      (src058[77] << 58) +
      (src058[78] << 58) +
      (src058[79] << 58) +
      (src058[80] << 58) +
      (src058[81] << 58) +
      (src058[82] << 58) +
      (src058[83] << 58) +
      (src058[84] << 58) +
      (src058[85] << 58) +
      (src058[86] << 58) +
      (src058[87] << 58) +
      (src058[88] << 58) +
      (src058[89] << 58) +
      (src058[90] << 58) +
      (src058[91] << 58) +
      (src058[92] << 58) +
      (src058[93] << 58) +
      (src058[94] << 58) +
      (src058[95] << 58) +
      (src058[96] << 58) +
      (src058[97] << 58) +
      (src058[98] << 58) +
      (src058[99] << 58) +
      (src058[100] << 58) +
      (src058[101] << 58) +
      (src058[102] << 58) +
      (src058[103] << 58) +
      (src058[104] << 58) +
      (src058[105] << 58) +
      (src058[106] << 58) +
      (src058[107] << 58) +
      (src058[108] << 58) +
      (src058[109] << 58) +
      (src058[110] << 58) +
      (src058[111] << 58) +
      (src058[112] << 58) +
      (src058[113] << 58) +
      (src058[114] << 58) +
      (src058[115] << 58) +
      (src058[116] << 58) +
      (src058[117] << 58) +
      (src058[118] << 58) +
      (src058[119] << 58) +
      (src058[120] << 58) +
      (src058[121] << 58) +
      (src058[122] << 58) +
      (src058[123] << 58) +
      (src058[124] << 58) +
      (src058[125] << 58) +
      (src058[126] << 58) +
      (src058[127] << 58) +
      (src059[0] << 59) +
      (src059[1] << 59) +
      (src059[2] << 59) +
      (src059[3] << 59) +
      (src059[4] << 59) +
      (src059[5] << 59) +
      (src059[6] << 59) +
      (src059[7] << 59) +
      (src059[8] << 59) +
      (src059[9] << 59) +
      (src059[10] << 59) +
      (src059[11] << 59) +
      (src059[12] << 59) +
      (src059[13] << 59) +
      (src059[14] << 59) +
      (src059[15] << 59) +
      (src059[16] << 59) +
      (src059[17] << 59) +
      (src059[18] << 59) +
      (src059[19] << 59) +
      (src059[20] << 59) +
      (src059[21] << 59) +
      (src059[22] << 59) +
      (src059[23] << 59) +
      (src059[24] << 59) +
      (src059[25] << 59) +
      (src059[26] << 59) +
      (src059[27] << 59) +
      (src059[28] << 59) +
      (src059[29] << 59) +
      (src059[30] << 59) +
      (src059[31] << 59) +
      (src059[32] << 59) +
      (src059[33] << 59) +
      (src059[34] << 59) +
      (src059[35] << 59) +
      (src059[36] << 59) +
      (src059[37] << 59) +
      (src059[38] << 59) +
      (src059[39] << 59) +
      (src059[40] << 59) +
      (src059[41] << 59) +
      (src059[42] << 59) +
      (src059[43] << 59) +
      (src059[44] << 59) +
      (src059[45] << 59) +
      (src059[46] << 59) +
      (src059[47] << 59) +
      (src059[48] << 59) +
      (src059[49] << 59) +
      (src059[50] << 59) +
      (src059[51] << 59) +
      (src059[52] << 59) +
      (src059[53] << 59) +
      (src059[54] << 59) +
      (src059[55] << 59) +
      (src059[56] << 59) +
      (src059[57] << 59) +
      (src059[58] << 59) +
      (src059[59] << 59) +
      (src059[60] << 59) +
      (src059[61] << 59) +
      (src059[62] << 59) +
      (src059[63] << 59) +
      (src059[64] << 59) +
      (src059[65] << 59) +
      (src059[66] << 59) +
      (src059[67] << 59) +
      (src059[68] << 59) +
      (src059[69] << 59) +
      (src059[70] << 59) +
      (src059[71] << 59) +
      (src059[72] << 59) +
      (src059[73] << 59) +
      (src059[74] << 59) +
      (src059[75] << 59) +
      (src059[76] << 59) +
      (src059[77] << 59) +
      (src059[78] << 59) +
      (src059[79] << 59) +
      (src059[80] << 59) +
      (src059[81] << 59) +
      (src059[82] << 59) +
      (src059[83] << 59) +
      (src059[84] << 59) +
      (src059[85] << 59) +
      (src059[86] << 59) +
      (src059[87] << 59) +
      (src059[88] << 59) +
      (src059[89] << 59) +
      (src059[90] << 59) +
      (src059[91] << 59) +
      (src059[92] << 59) +
      (src059[93] << 59) +
      (src059[94] << 59) +
      (src059[95] << 59) +
      (src059[96] << 59) +
      (src059[97] << 59) +
      (src059[98] << 59) +
      (src059[99] << 59) +
      (src059[100] << 59) +
      (src059[101] << 59) +
      (src059[102] << 59) +
      (src059[103] << 59) +
      (src059[104] << 59) +
      (src059[105] << 59) +
      (src059[106] << 59) +
      (src059[107] << 59) +
      (src059[108] << 59) +
      (src059[109] << 59) +
      (src059[110] << 59) +
      (src059[111] << 59) +
      (src059[112] << 59) +
      (src059[113] << 59) +
      (src059[114] << 59) +
      (src059[115] << 59) +
      (src059[116] << 59) +
      (src059[117] << 59) +
      (src059[118] << 59) +
      (src059[119] << 59) +
      (src059[120] << 59) +
      (src059[121] << 59) +
      (src059[122] << 59) +
      (src059[123] << 59) +
      (src059[124] << 59) +
      (src059[125] << 59) +
      (src059[126] << 59) +
      (src059[127] << 59) +
      (src060[0] << 60) +
      (src060[1] << 60) +
      (src060[2] << 60) +
      (src060[3] << 60) +
      (src060[4] << 60) +
      (src060[5] << 60) +
      (src060[6] << 60) +
      (src060[7] << 60) +
      (src060[8] << 60) +
      (src060[9] << 60) +
      (src060[10] << 60) +
      (src060[11] << 60) +
      (src060[12] << 60) +
      (src060[13] << 60) +
      (src060[14] << 60) +
      (src060[15] << 60) +
      (src060[16] << 60) +
      (src060[17] << 60) +
      (src060[18] << 60) +
      (src060[19] << 60) +
      (src060[20] << 60) +
      (src060[21] << 60) +
      (src060[22] << 60) +
      (src060[23] << 60) +
      (src060[24] << 60) +
      (src060[25] << 60) +
      (src060[26] << 60) +
      (src060[27] << 60) +
      (src060[28] << 60) +
      (src060[29] << 60) +
      (src060[30] << 60) +
      (src060[31] << 60) +
      (src060[32] << 60) +
      (src060[33] << 60) +
      (src060[34] << 60) +
      (src060[35] << 60) +
      (src060[36] << 60) +
      (src060[37] << 60) +
      (src060[38] << 60) +
      (src060[39] << 60) +
      (src060[40] << 60) +
      (src060[41] << 60) +
      (src060[42] << 60) +
      (src060[43] << 60) +
      (src060[44] << 60) +
      (src060[45] << 60) +
      (src060[46] << 60) +
      (src060[47] << 60) +
      (src060[48] << 60) +
      (src060[49] << 60) +
      (src060[50] << 60) +
      (src060[51] << 60) +
      (src060[52] << 60) +
      (src060[53] << 60) +
      (src060[54] << 60) +
      (src060[55] << 60) +
      (src060[56] << 60) +
      (src060[57] << 60) +
      (src060[58] << 60) +
      (src060[59] << 60) +
      (src060[60] << 60) +
      (src060[61] << 60) +
      (src060[62] << 60) +
      (src060[63] << 60) +
      (src060[64] << 60) +
      (src060[65] << 60) +
      (src060[66] << 60) +
      (src060[67] << 60) +
      (src060[68] << 60) +
      (src060[69] << 60) +
      (src060[70] << 60) +
      (src060[71] << 60) +
      (src060[72] << 60) +
      (src060[73] << 60) +
      (src060[74] << 60) +
      (src060[75] << 60) +
      (src060[76] << 60) +
      (src060[77] << 60) +
      (src060[78] << 60) +
      (src060[79] << 60) +
      (src060[80] << 60) +
      (src060[81] << 60) +
      (src060[82] << 60) +
      (src060[83] << 60) +
      (src060[84] << 60) +
      (src060[85] << 60) +
      (src060[86] << 60) +
      (src060[87] << 60) +
      (src060[88] << 60) +
      (src060[89] << 60) +
      (src060[90] << 60) +
      (src060[91] << 60) +
      (src060[92] << 60) +
      (src060[93] << 60) +
      (src060[94] << 60) +
      (src060[95] << 60) +
      (src060[96] << 60) +
      (src060[97] << 60) +
      (src060[98] << 60) +
      (src060[99] << 60) +
      (src060[100] << 60) +
      (src060[101] << 60) +
      (src060[102] << 60) +
      (src060[103] << 60) +
      (src060[104] << 60) +
      (src060[105] << 60) +
      (src060[106] << 60) +
      (src060[107] << 60) +
      (src060[108] << 60) +
      (src060[109] << 60) +
      (src060[110] << 60) +
      (src060[111] << 60) +
      (src060[112] << 60) +
      (src060[113] << 60) +
      (src060[114] << 60) +
      (src060[115] << 60) +
      (src060[116] << 60) +
      (src060[117] << 60) +
      (src060[118] << 60) +
      (src060[119] << 60) +
      (src060[120] << 60) +
      (src060[121] << 60) +
      (src060[122] << 60) +
      (src060[123] << 60) +
      (src060[124] << 60) +
      (src060[125] << 60) +
      (src060[126] << 60) +
      (src060[127] << 60) +
      (src061[0] << 61) +
      (src061[1] << 61) +
      (src061[2] << 61) +
      (src061[3] << 61) +
      (src061[4] << 61) +
      (src061[5] << 61) +
      (src061[6] << 61) +
      (src061[7] << 61) +
      (src061[8] << 61) +
      (src061[9] << 61) +
      (src061[10] << 61) +
      (src061[11] << 61) +
      (src061[12] << 61) +
      (src061[13] << 61) +
      (src061[14] << 61) +
      (src061[15] << 61) +
      (src061[16] << 61) +
      (src061[17] << 61) +
      (src061[18] << 61) +
      (src061[19] << 61) +
      (src061[20] << 61) +
      (src061[21] << 61) +
      (src061[22] << 61) +
      (src061[23] << 61) +
      (src061[24] << 61) +
      (src061[25] << 61) +
      (src061[26] << 61) +
      (src061[27] << 61) +
      (src061[28] << 61) +
      (src061[29] << 61) +
      (src061[30] << 61) +
      (src061[31] << 61) +
      (src061[32] << 61) +
      (src061[33] << 61) +
      (src061[34] << 61) +
      (src061[35] << 61) +
      (src061[36] << 61) +
      (src061[37] << 61) +
      (src061[38] << 61) +
      (src061[39] << 61) +
      (src061[40] << 61) +
      (src061[41] << 61) +
      (src061[42] << 61) +
      (src061[43] << 61) +
      (src061[44] << 61) +
      (src061[45] << 61) +
      (src061[46] << 61) +
      (src061[47] << 61) +
      (src061[48] << 61) +
      (src061[49] << 61) +
      (src061[50] << 61) +
      (src061[51] << 61) +
      (src061[52] << 61) +
      (src061[53] << 61) +
      (src061[54] << 61) +
      (src061[55] << 61) +
      (src061[56] << 61) +
      (src061[57] << 61) +
      (src061[58] << 61) +
      (src061[59] << 61) +
      (src061[60] << 61) +
      (src061[61] << 61) +
      (src061[62] << 61) +
      (src061[63] << 61) +
      (src061[64] << 61) +
      (src061[65] << 61) +
      (src061[66] << 61) +
      (src061[67] << 61) +
      (src061[68] << 61) +
      (src061[69] << 61) +
      (src061[70] << 61) +
      (src061[71] << 61) +
      (src061[72] << 61) +
      (src061[73] << 61) +
      (src061[74] << 61) +
      (src061[75] << 61) +
      (src061[76] << 61) +
      (src061[77] << 61) +
      (src061[78] << 61) +
      (src061[79] << 61) +
      (src061[80] << 61) +
      (src061[81] << 61) +
      (src061[82] << 61) +
      (src061[83] << 61) +
      (src061[84] << 61) +
      (src061[85] << 61) +
      (src061[86] << 61) +
      (src061[87] << 61) +
      (src061[88] << 61) +
      (src061[89] << 61) +
      (src061[90] << 61) +
      (src061[91] << 61) +
      (src061[92] << 61) +
      (src061[93] << 61) +
      (src061[94] << 61) +
      (src061[95] << 61) +
      (src061[96] << 61) +
      (src061[97] << 61) +
      (src061[98] << 61) +
      (src061[99] << 61) +
      (src061[100] << 61) +
      (src061[101] << 61) +
      (src061[102] << 61) +
      (src061[103] << 61) +
      (src061[104] << 61) +
      (src061[105] << 61) +
      (src061[106] << 61) +
      (src061[107] << 61) +
      (src061[108] << 61) +
      (src061[109] << 61) +
      (src061[110] << 61) +
      (src061[111] << 61) +
      (src061[112] << 61) +
      (src061[113] << 61) +
      (src061[114] << 61) +
      (src061[115] << 61) +
      (src061[116] << 61) +
      (src061[117] << 61) +
      (src061[118] << 61) +
      (src061[119] << 61) +
      (src061[120] << 61) +
      (src061[121] << 61) +
      (src061[122] << 61) +
      (src061[123] << 61) +
      (src061[124] << 61) +
      (src061[125] << 61) +
      (src061[126] << 61) +
      (src061[127] << 61) +
      (src062[0] << 62) +
      (src062[1] << 62) +
      (src062[2] << 62) +
      (src062[3] << 62) +
      (src062[4] << 62) +
      (src062[5] << 62) +
      (src062[6] << 62) +
      (src062[7] << 62) +
      (src062[8] << 62) +
      (src062[9] << 62) +
      (src062[10] << 62) +
      (src062[11] << 62) +
      (src062[12] << 62) +
      (src062[13] << 62) +
      (src062[14] << 62) +
      (src062[15] << 62) +
      (src062[16] << 62) +
      (src062[17] << 62) +
      (src062[18] << 62) +
      (src062[19] << 62) +
      (src062[20] << 62) +
      (src062[21] << 62) +
      (src062[22] << 62) +
      (src062[23] << 62) +
      (src062[24] << 62) +
      (src062[25] << 62) +
      (src062[26] << 62) +
      (src062[27] << 62) +
      (src062[28] << 62) +
      (src062[29] << 62) +
      (src062[30] << 62) +
      (src062[31] << 62) +
      (src062[32] << 62) +
      (src062[33] << 62) +
      (src062[34] << 62) +
      (src062[35] << 62) +
      (src062[36] << 62) +
      (src062[37] << 62) +
      (src062[38] << 62) +
      (src062[39] << 62) +
      (src062[40] << 62) +
      (src062[41] << 62) +
      (src062[42] << 62) +
      (src062[43] << 62) +
      (src062[44] << 62) +
      (src062[45] << 62) +
      (src062[46] << 62) +
      (src062[47] << 62) +
      (src062[48] << 62) +
      (src062[49] << 62) +
      (src062[50] << 62) +
      (src062[51] << 62) +
      (src062[52] << 62) +
      (src062[53] << 62) +
      (src062[54] << 62) +
      (src062[55] << 62) +
      (src062[56] << 62) +
      (src062[57] << 62) +
      (src062[58] << 62) +
      (src062[59] << 62) +
      (src062[60] << 62) +
      (src062[61] << 62) +
      (src062[62] << 62) +
      (src062[63] << 62) +
      (src062[64] << 62) +
      (src062[65] << 62) +
      (src062[66] << 62) +
      (src062[67] << 62) +
      (src062[68] << 62) +
      (src062[69] << 62) +
      (src062[70] << 62) +
      (src062[71] << 62) +
      (src062[72] << 62) +
      (src062[73] << 62) +
      (src062[74] << 62) +
      (src062[75] << 62) +
      (src062[76] << 62) +
      (src062[77] << 62) +
      (src062[78] << 62) +
      (src062[79] << 62) +
      (src062[80] << 62) +
      (src062[81] << 62) +
      (src062[82] << 62) +
      (src062[83] << 62) +
      (src062[84] << 62) +
      (src062[85] << 62) +
      (src062[86] << 62) +
      (src062[87] << 62) +
      (src062[88] << 62) +
      (src062[89] << 62) +
      (src062[90] << 62) +
      (src062[91] << 62) +
      (src062[92] << 62) +
      (src062[93] << 62) +
      (src062[94] << 62) +
      (src062[95] << 62) +
      (src062[96] << 62) +
      (src062[97] << 62) +
      (src062[98] << 62) +
      (src062[99] << 62) +
      (src062[100] << 62) +
      (src062[101] << 62) +
      (src062[102] << 62) +
      (src062[103] << 62) +
      (src062[104] << 62) +
      (src062[105] << 62) +
      (src062[106] << 62) +
      (src062[107] << 62) +
      (src062[108] << 62) +
      (src062[109] << 62) +
      (src062[110] << 62) +
      (src062[111] << 62) +
      (src062[112] << 62) +
      (src062[113] << 62) +
      (src062[114] << 62) +
      (src062[115] << 62) +
      (src062[116] << 62) +
      (src062[117] << 62) +
      (src062[118] << 62) +
      (src062[119] << 62) +
      (src062[120] << 62) +
      (src062[121] << 62) +
      (src062[122] << 62) +
      (src062[123] << 62) +
      (src062[124] << 62) +
      (src062[125] << 62) +
      (src062[126] << 62) +
      (src062[127] << 62) +
      (src063[0] << 63) +
      (src063[1] << 63) +
      (src063[2] << 63) +
      (src063[3] << 63) +
      (src063[4] << 63) +
      (src063[5] << 63) +
      (src063[6] << 63) +
      (src063[7] << 63) +
      (src063[8] << 63) +
      (src063[9] << 63) +
      (src063[10] << 63) +
      (src063[11] << 63) +
      (src063[12] << 63) +
      (src063[13] << 63) +
      (src063[14] << 63) +
      (src063[15] << 63) +
      (src063[16] << 63) +
      (src063[17] << 63) +
      (src063[18] << 63) +
      (src063[19] << 63) +
      (src063[20] << 63) +
      (src063[21] << 63) +
      (src063[22] << 63) +
      (src063[23] << 63) +
      (src063[24] << 63) +
      (src063[25] << 63) +
      (src063[26] << 63) +
      (src063[27] << 63) +
      (src063[28] << 63) +
      (src063[29] << 63) +
      (src063[30] << 63) +
      (src063[31] << 63) +
      (src063[32] << 63) +
      (src063[33] << 63) +
      (src063[34] << 63) +
      (src063[35] << 63) +
      (src063[36] << 63) +
      (src063[37] << 63) +
      (src063[38] << 63) +
      (src063[39] << 63) +
      (src063[40] << 63) +
      (src063[41] << 63) +
      (src063[42] << 63) +
      (src063[43] << 63) +
      (src063[44] << 63) +
      (src063[45] << 63) +
      (src063[46] << 63) +
      (src063[47] << 63) +
      (src063[48] << 63) +
      (src063[49] << 63) +
      (src063[50] << 63) +
      (src063[51] << 63) +
      (src063[52] << 63) +
      (src063[53] << 63) +
      (src063[54] << 63) +
      (src063[55] << 63) +
      (src063[56] << 63) +
      (src063[57] << 63) +
      (src063[58] << 63) +
      (src063[59] << 63) +
      (src063[60] << 63) +
      (src063[61] << 63) +
      (src063[62] << 63) +
      (src063[63] << 63) +
      (src063[64] << 63) +
      (src063[65] << 63) +
      (src063[66] << 63) +
      (src063[67] << 63) +
      (src063[68] << 63) +
      (src063[69] << 63) +
      (src063[70] << 63) +
      (src063[71] << 63) +
      (src063[72] << 63) +
      (src063[73] << 63) +
      (src063[74] << 63) +
      (src063[75] << 63) +
      (src063[76] << 63) +
      (src063[77] << 63) +
      (src063[78] << 63) +
      (src063[79] << 63) +
      (src063[80] << 63) +
      (src063[81] << 63) +
      (src063[82] << 63) +
      (src063[83] << 63) +
      (src063[84] << 63) +
      (src063[85] << 63) +
      (src063[86] << 63) +
      (src063[87] << 63) +
      (src063[88] << 63) +
      (src063[89] << 63) +
      (src063[90] << 63) +
      (src063[91] << 63) +
      (src063[92] << 63) +
      (src063[93] << 63) +
      (src063[94] << 63) +
      (src063[95] << 63) +
      (src063[96] << 63) +
      (src063[97] << 63) +
      (src063[98] << 63) +
      (src063[99] << 63) +
      (src063[100] << 63) +
      (src063[101] << 63) +
      (src063[102] << 63) +
      (src063[103] << 63) +
      (src063[104] << 63) +
      (src063[105] << 63) +
      (src063[106] << 63) +
      (src063[107] << 63) +
      (src063[108] << 63) +
      (src063[109] << 63) +
      (src063[110] << 63) +
      (src063[111] << 63) +
      (src063[112] << 63) +
      (src063[113] << 63) +
      (src063[114] << 63) +
      (src063[115] << 63) +
      (src063[116] << 63) +
      (src063[117] << 63) +
      (src063[118] << 63) +
      (src063[119] << 63) +
      (src063[120] << 63) +
      (src063[121] << 63) +
      (src063[122] << 63) +
      (src063[123] << 63) +
      (src063[124] << 63) +
      (src063[125] << 63) +
      (src063[126] << 63) +
      (src063[127] << 63) +
      (src064[0] << 64) +
      (src064[1] << 64) +
      (src064[2] << 64) +
      (src064[3] << 64) +
      (src064[4] << 64) +
      (src064[5] << 64) +
      (src064[6] << 64) +
      (src064[7] << 64) +
      (src064[8] << 64) +
      (src064[9] << 64) +
      (src064[10] << 64) +
      (src064[11] << 64) +
      (src064[12] << 64) +
      (src064[13] << 64) +
      (src064[14] << 64) +
      (src064[15] << 64) +
      (src064[16] << 64) +
      (src064[17] << 64) +
      (src064[18] << 64) +
      (src064[19] << 64) +
      (src064[20] << 64) +
      (src064[21] << 64) +
      (src064[22] << 64) +
      (src064[23] << 64) +
      (src064[24] << 64) +
      (src064[25] << 64) +
      (src064[26] << 64) +
      (src064[27] << 64) +
      (src064[28] << 64) +
      (src064[29] << 64) +
      (src064[30] << 64) +
      (src064[31] << 64) +
      (src064[32] << 64) +
      (src064[33] << 64) +
      (src064[34] << 64) +
      (src064[35] << 64) +
      (src064[36] << 64) +
      (src064[37] << 64) +
      (src064[38] << 64) +
      (src064[39] << 64) +
      (src064[40] << 64) +
      (src064[41] << 64) +
      (src064[42] << 64) +
      (src064[43] << 64) +
      (src064[44] << 64) +
      (src064[45] << 64) +
      (src064[46] << 64) +
      (src064[47] << 64) +
      (src064[48] << 64) +
      (src064[49] << 64) +
      (src064[50] << 64) +
      (src064[51] << 64) +
      (src064[52] << 64) +
      (src064[53] << 64) +
      (src064[54] << 64) +
      (src064[55] << 64) +
      (src064[56] << 64) +
      (src064[57] << 64) +
      (src064[58] << 64) +
      (src064[59] << 64) +
      (src064[60] << 64) +
      (src064[61] << 64) +
      (src064[62] << 64) +
      (src064[63] << 64) +
      (src064[64] << 64) +
      (src064[65] << 64) +
      (src064[66] << 64) +
      (src064[67] << 64) +
      (src064[68] << 64) +
      (src064[69] << 64) +
      (src064[70] << 64) +
      (src064[71] << 64) +
      (src064[72] << 64) +
      (src064[73] << 64) +
      (src064[74] << 64) +
      (src064[75] << 64) +
      (src064[76] << 64) +
      (src064[77] << 64) +
      (src064[78] << 64) +
      (src064[79] << 64) +
      (src064[80] << 64) +
      (src064[81] << 64) +
      (src064[82] << 64) +
      (src064[83] << 64) +
      (src064[84] << 64) +
      (src064[85] << 64) +
      (src064[86] << 64) +
      (src064[87] << 64) +
      (src064[88] << 64) +
      (src064[89] << 64) +
      (src064[90] << 64) +
      (src064[91] << 64) +
      (src064[92] << 64) +
      (src064[93] << 64) +
      (src064[94] << 64) +
      (src064[95] << 64) +
      (src064[96] << 64) +
      (src064[97] << 64) +
      (src064[98] << 64) +
      (src064[99] << 64) +
      (src064[100] << 64) +
      (src064[101] << 64) +
      (src064[102] << 64) +
      (src064[103] << 64) +
      (src064[104] << 64) +
      (src064[105] << 64) +
      (src064[106] << 64) +
      (src064[107] << 64) +
      (src064[108] << 64) +
      (src064[109] << 64) +
      (src064[110] << 64) +
      (src064[111] << 64) +
      (src064[112] << 64) +
      (src064[113] << 64) +
      (src064[114] << 64) +
      (src064[115] << 64) +
      (src064[116] << 64) +
      (src064[117] << 64) +
      (src064[118] << 64) +
      (src064[119] << 64) +
      (src064[120] << 64) +
      (src064[121] << 64) +
      (src064[122] << 64) +
      (src064[123] << 64) +
      (src064[124] << 64) +
      (src064[125] << 64) +
      (src064[126] << 64) +
      (src064[127] << 64) +
      (src065[0] << 65) +
      (src065[1] << 65) +
      (src065[2] << 65) +
      (src065[3] << 65) +
      (src065[4] << 65) +
      (src065[5] << 65) +
      (src065[6] << 65) +
      (src065[7] << 65) +
      (src065[8] << 65) +
      (src065[9] << 65) +
      (src065[10] << 65) +
      (src065[11] << 65) +
      (src065[12] << 65) +
      (src065[13] << 65) +
      (src065[14] << 65) +
      (src065[15] << 65) +
      (src065[16] << 65) +
      (src065[17] << 65) +
      (src065[18] << 65) +
      (src065[19] << 65) +
      (src065[20] << 65) +
      (src065[21] << 65) +
      (src065[22] << 65) +
      (src065[23] << 65) +
      (src065[24] << 65) +
      (src065[25] << 65) +
      (src065[26] << 65) +
      (src065[27] << 65) +
      (src065[28] << 65) +
      (src065[29] << 65) +
      (src065[30] << 65) +
      (src065[31] << 65) +
      (src065[32] << 65) +
      (src065[33] << 65) +
      (src065[34] << 65) +
      (src065[35] << 65) +
      (src065[36] << 65) +
      (src065[37] << 65) +
      (src065[38] << 65) +
      (src065[39] << 65) +
      (src065[40] << 65) +
      (src065[41] << 65) +
      (src065[42] << 65) +
      (src065[43] << 65) +
      (src065[44] << 65) +
      (src065[45] << 65) +
      (src065[46] << 65) +
      (src065[47] << 65) +
      (src065[48] << 65) +
      (src065[49] << 65) +
      (src065[50] << 65) +
      (src065[51] << 65) +
      (src065[52] << 65) +
      (src065[53] << 65) +
      (src065[54] << 65) +
      (src065[55] << 65) +
      (src065[56] << 65) +
      (src065[57] << 65) +
      (src065[58] << 65) +
      (src065[59] << 65) +
      (src065[60] << 65) +
      (src065[61] << 65) +
      (src065[62] << 65) +
      (src065[63] << 65) +
      (src065[64] << 65) +
      (src065[65] << 65) +
      (src065[66] << 65) +
      (src065[67] << 65) +
      (src065[68] << 65) +
      (src065[69] << 65) +
      (src065[70] << 65) +
      (src065[71] << 65) +
      (src065[72] << 65) +
      (src065[73] << 65) +
      (src065[74] << 65) +
      (src065[75] << 65) +
      (src065[76] << 65) +
      (src065[77] << 65) +
      (src065[78] << 65) +
      (src065[79] << 65) +
      (src065[80] << 65) +
      (src065[81] << 65) +
      (src065[82] << 65) +
      (src065[83] << 65) +
      (src065[84] << 65) +
      (src065[85] << 65) +
      (src065[86] << 65) +
      (src065[87] << 65) +
      (src065[88] << 65) +
      (src065[89] << 65) +
      (src065[90] << 65) +
      (src065[91] << 65) +
      (src065[92] << 65) +
      (src065[93] << 65) +
      (src065[94] << 65) +
      (src065[95] << 65) +
      (src065[96] << 65) +
      (src065[97] << 65) +
      (src065[98] << 65) +
      (src065[99] << 65) +
      (src065[100] << 65) +
      (src065[101] << 65) +
      (src065[102] << 65) +
      (src065[103] << 65) +
      (src065[104] << 65) +
      (src065[105] << 65) +
      (src065[106] << 65) +
      (src065[107] << 65) +
      (src065[108] << 65) +
      (src065[109] << 65) +
      (src065[110] << 65) +
      (src065[111] << 65) +
      (src065[112] << 65) +
      (src065[113] << 65) +
      (src065[114] << 65) +
      (src065[115] << 65) +
      (src065[116] << 65) +
      (src065[117] << 65) +
      (src065[118] << 65) +
      (src065[119] << 65) +
      (src065[120] << 65) +
      (src065[121] << 65) +
      (src065[122] << 65) +
      (src065[123] << 65) +
      (src065[124] << 65) +
      (src065[125] << 65) +
      (src065[126] << 65) +
      (src065[127] << 65) +
      (src066[0] << 66) +
      (src066[1] << 66) +
      (src066[2] << 66) +
      (src066[3] << 66) +
      (src066[4] << 66) +
      (src066[5] << 66) +
      (src066[6] << 66) +
      (src066[7] << 66) +
      (src066[8] << 66) +
      (src066[9] << 66) +
      (src066[10] << 66) +
      (src066[11] << 66) +
      (src066[12] << 66) +
      (src066[13] << 66) +
      (src066[14] << 66) +
      (src066[15] << 66) +
      (src066[16] << 66) +
      (src066[17] << 66) +
      (src066[18] << 66) +
      (src066[19] << 66) +
      (src066[20] << 66) +
      (src066[21] << 66) +
      (src066[22] << 66) +
      (src066[23] << 66) +
      (src066[24] << 66) +
      (src066[25] << 66) +
      (src066[26] << 66) +
      (src066[27] << 66) +
      (src066[28] << 66) +
      (src066[29] << 66) +
      (src066[30] << 66) +
      (src066[31] << 66) +
      (src066[32] << 66) +
      (src066[33] << 66) +
      (src066[34] << 66) +
      (src066[35] << 66) +
      (src066[36] << 66) +
      (src066[37] << 66) +
      (src066[38] << 66) +
      (src066[39] << 66) +
      (src066[40] << 66) +
      (src066[41] << 66) +
      (src066[42] << 66) +
      (src066[43] << 66) +
      (src066[44] << 66) +
      (src066[45] << 66) +
      (src066[46] << 66) +
      (src066[47] << 66) +
      (src066[48] << 66) +
      (src066[49] << 66) +
      (src066[50] << 66) +
      (src066[51] << 66) +
      (src066[52] << 66) +
      (src066[53] << 66) +
      (src066[54] << 66) +
      (src066[55] << 66) +
      (src066[56] << 66) +
      (src066[57] << 66) +
      (src066[58] << 66) +
      (src066[59] << 66) +
      (src066[60] << 66) +
      (src066[61] << 66) +
      (src066[62] << 66) +
      (src066[63] << 66) +
      (src066[64] << 66) +
      (src066[65] << 66) +
      (src066[66] << 66) +
      (src066[67] << 66) +
      (src066[68] << 66) +
      (src066[69] << 66) +
      (src066[70] << 66) +
      (src066[71] << 66) +
      (src066[72] << 66) +
      (src066[73] << 66) +
      (src066[74] << 66) +
      (src066[75] << 66) +
      (src066[76] << 66) +
      (src066[77] << 66) +
      (src066[78] << 66) +
      (src066[79] << 66) +
      (src066[80] << 66) +
      (src066[81] << 66) +
      (src066[82] << 66) +
      (src066[83] << 66) +
      (src066[84] << 66) +
      (src066[85] << 66) +
      (src066[86] << 66) +
      (src066[87] << 66) +
      (src066[88] << 66) +
      (src066[89] << 66) +
      (src066[90] << 66) +
      (src066[91] << 66) +
      (src066[92] << 66) +
      (src066[93] << 66) +
      (src066[94] << 66) +
      (src066[95] << 66) +
      (src066[96] << 66) +
      (src066[97] << 66) +
      (src066[98] << 66) +
      (src066[99] << 66) +
      (src066[100] << 66) +
      (src066[101] << 66) +
      (src066[102] << 66) +
      (src066[103] << 66) +
      (src066[104] << 66) +
      (src066[105] << 66) +
      (src066[106] << 66) +
      (src066[107] << 66) +
      (src066[108] << 66) +
      (src066[109] << 66) +
      (src066[110] << 66) +
      (src066[111] << 66) +
      (src066[112] << 66) +
      (src066[113] << 66) +
      (src066[114] << 66) +
      (src066[115] << 66) +
      (src066[116] << 66) +
      (src066[117] << 66) +
      (src066[118] << 66) +
      (src066[119] << 66) +
      (src066[120] << 66) +
      (src066[121] << 66) +
      (src066[122] << 66) +
      (src066[123] << 66) +
      (src066[124] << 66) +
      (src066[125] << 66) +
      (src066[126] << 66) +
      (src066[127] << 66) +
      (src067[0] << 67) +
      (src067[1] << 67) +
      (src067[2] << 67) +
      (src067[3] << 67) +
      (src067[4] << 67) +
      (src067[5] << 67) +
      (src067[6] << 67) +
      (src067[7] << 67) +
      (src067[8] << 67) +
      (src067[9] << 67) +
      (src067[10] << 67) +
      (src067[11] << 67) +
      (src067[12] << 67) +
      (src067[13] << 67) +
      (src067[14] << 67) +
      (src067[15] << 67) +
      (src067[16] << 67) +
      (src067[17] << 67) +
      (src067[18] << 67) +
      (src067[19] << 67) +
      (src067[20] << 67) +
      (src067[21] << 67) +
      (src067[22] << 67) +
      (src067[23] << 67) +
      (src067[24] << 67) +
      (src067[25] << 67) +
      (src067[26] << 67) +
      (src067[27] << 67) +
      (src067[28] << 67) +
      (src067[29] << 67) +
      (src067[30] << 67) +
      (src067[31] << 67) +
      (src067[32] << 67) +
      (src067[33] << 67) +
      (src067[34] << 67) +
      (src067[35] << 67) +
      (src067[36] << 67) +
      (src067[37] << 67) +
      (src067[38] << 67) +
      (src067[39] << 67) +
      (src067[40] << 67) +
      (src067[41] << 67) +
      (src067[42] << 67) +
      (src067[43] << 67) +
      (src067[44] << 67) +
      (src067[45] << 67) +
      (src067[46] << 67) +
      (src067[47] << 67) +
      (src067[48] << 67) +
      (src067[49] << 67) +
      (src067[50] << 67) +
      (src067[51] << 67) +
      (src067[52] << 67) +
      (src067[53] << 67) +
      (src067[54] << 67) +
      (src067[55] << 67) +
      (src067[56] << 67) +
      (src067[57] << 67) +
      (src067[58] << 67) +
      (src067[59] << 67) +
      (src067[60] << 67) +
      (src067[61] << 67) +
      (src067[62] << 67) +
      (src067[63] << 67) +
      (src067[64] << 67) +
      (src067[65] << 67) +
      (src067[66] << 67) +
      (src067[67] << 67) +
      (src067[68] << 67) +
      (src067[69] << 67) +
      (src067[70] << 67) +
      (src067[71] << 67) +
      (src067[72] << 67) +
      (src067[73] << 67) +
      (src067[74] << 67) +
      (src067[75] << 67) +
      (src067[76] << 67) +
      (src067[77] << 67) +
      (src067[78] << 67) +
      (src067[79] << 67) +
      (src067[80] << 67) +
      (src067[81] << 67) +
      (src067[82] << 67) +
      (src067[83] << 67) +
      (src067[84] << 67) +
      (src067[85] << 67) +
      (src067[86] << 67) +
      (src067[87] << 67) +
      (src067[88] << 67) +
      (src067[89] << 67) +
      (src067[90] << 67) +
      (src067[91] << 67) +
      (src067[92] << 67) +
      (src067[93] << 67) +
      (src067[94] << 67) +
      (src067[95] << 67) +
      (src067[96] << 67) +
      (src067[97] << 67) +
      (src067[98] << 67) +
      (src067[99] << 67) +
      (src067[100] << 67) +
      (src067[101] << 67) +
      (src067[102] << 67) +
      (src067[103] << 67) +
      (src067[104] << 67) +
      (src067[105] << 67) +
      (src067[106] << 67) +
      (src067[107] << 67) +
      (src067[108] << 67) +
      (src067[109] << 67) +
      (src067[110] << 67) +
      (src067[111] << 67) +
      (src067[112] << 67) +
      (src067[113] << 67) +
      (src067[114] << 67) +
      (src067[115] << 67) +
      (src067[116] << 67) +
      (src067[117] << 67) +
      (src067[118] << 67) +
      (src067[119] << 67) +
      (src067[120] << 67) +
      (src067[121] << 67) +
      (src067[122] << 67) +
      (src067[123] << 67) +
      (src067[124] << 67) +
      (src067[125] << 67) +
      (src067[126] << 67) +
      (src067[127] << 67) +
      (src068[0] << 68) +
      (src068[1] << 68) +
      (src068[2] << 68) +
      (src068[3] << 68) +
      (src068[4] << 68) +
      (src068[5] << 68) +
      (src068[6] << 68) +
      (src068[7] << 68) +
      (src068[8] << 68) +
      (src068[9] << 68) +
      (src068[10] << 68) +
      (src068[11] << 68) +
      (src068[12] << 68) +
      (src068[13] << 68) +
      (src068[14] << 68) +
      (src068[15] << 68) +
      (src068[16] << 68) +
      (src068[17] << 68) +
      (src068[18] << 68) +
      (src068[19] << 68) +
      (src068[20] << 68) +
      (src068[21] << 68) +
      (src068[22] << 68) +
      (src068[23] << 68) +
      (src068[24] << 68) +
      (src068[25] << 68) +
      (src068[26] << 68) +
      (src068[27] << 68) +
      (src068[28] << 68) +
      (src068[29] << 68) +
      (src068[30] << 68) +
      (src068[31] << 68) +
      (src068[32] << 68) +
      (src068[33] << 68) +
      (src068[34] << 68) +
      (src068[35] << 68) +
      (src068[36] << 68) +
      (src068[37] << 68) +
      (src068[38] << 68) +
      (src068[39] << 68) +
      (src068[40] << 68) +
      (src068[41] << 68) +
      (src068[42] << 68) +
      (src068[43] << 68) +
      (src068[44] << 68) +
      (src068[45] << 68) +
      (src068[46] << 68) +
      (src068[47] << 68) +
      (src068[48] << 68) +
      (src068[49] << 68) +
      (src068[50] << 68) +
      (src068[51] << 68) +
      (src068[52] << 68) +
      (src068[53] << 68) +
      (src068[54] << 68) +
      (src068[55] << 68) +
      (src068[56] << 68) +
      (src068[57] << 68) +
      (src068[58] << 68) +
      (src068[59] << 68) +
      (src068[60] << 68) +
      (src068[61] << 68) +
      (src068[62] << 68) +
      (src068[63] << 68) +
      (src068[64] << 68) +
      (src068[65] << 68) +
      (src068[66] << 68) +
      (src068[67] << 68) +
      (src068[68] << 68) +
      (src068[69] << 68) +
      (src068[70] << 68) +
      (src068[71] << 68) +
      (src068[72] << 68) +
      (src068[73] << 68) +
      (src068[74] << 68) +
      (src068[75] << 68) +
      (src068[76] << 68) +
      (src068[77] << 68) +
      (src068[78] << 68) +
      (src068[79] << 68) +
      (src068[80] << 68) +
      (src068[81] << 68) +
      (src068[82] << 68) +
      (src068[83] << 68) +
      (src068[84] << 68) +
      (src068[85] << 68) +
      (src068[86] << 68) +
      (src068[87] << 68) +
      (src068[88] << 68) +
      (src068[89] << 68) +
      (src068[90] << 68) +
      (src068[91] << 68) +
      (src068[92] << 68) +
      (src068[93] << 68) +
      (src068[94] << 68) +
      (src068[95] << 68) +
      (src068[96] << 68) +
      (src068[97] << 68) +
      (src068[98] << 68) +
      (src068[99] << 68) +
      (src068[100] << 68) +
      (src068[101] << 68) +
      (src068[102] << 68) +
      (src068[103] << 68) +
      (src068[104] << 68) +
      (src068[105] << 68) +
      (src068[106] << 68) +
      (src068[107] << 68) +
      (src068[108] << 68) +
      (src068[109] << 68) +
      (src068[110] << 68) +
      (src068[111] << 68) +
      (src068[112] << 68) +
      (src068[113] << 68) +
      (src068[114] << 68) +
      (src068[115] << 68) +
      (src068[116] << 68) +
      (src068[117] << 68) +
      (src068[118] << 68) +
      (src068[119] << 68) +
      (src068[120] << 68) +
      (src068[121] << 68) +
      (src068[122] << 68) +
      (src068[123] << 68) +
      (src068[124] << 68) +
      (src068[125] << 68) +
      (src068[126] << 68) +
      (src068[127] << 68) +
      (src069[0] << 69) +
      (src069[1] << 69) +
      (src069[2] << 69) +
      (src069[3] << 69) +
      (src069[4] << 69) +
      (src069[5] << 69) +
      (src069[6] << 69) +
      (src069[7] << 69) +
      (src069[8] << 69) +
      (src069[9] << 69) +
      (src069[10] << 69) +
      (src069[11] << 69) +
      (src069[12] << 69) +
      (src069[13] << 69) +
      (src069[14] << 69) +
      (src069[15] << 69) +
      (src069[16] << 69) +
      (src069[17] << 69) +
      (src069[18] << 69) +
      (src069[19] << 69) +
      (src069[20] << 69) +
      (src069[21] << 69) +
      (src069[22] << 69) +
      (src069[23] << 69) +
      (src069[24] << 69) +
      (src069[25] << 69) +
      (src069[26] << 69) +
      (src069[27] << 69) +
      (src069[28] << 69) +
      (src069[29] << 69) +
      (src069[30] << 69) +
      (src069[31] << 69) +
      (src069[32] << 69) +
      (src069[33] << 69) +
      (src069[34] << 69) +
      (src069[35] << 69) +
      (src069[36] << 69) +
      (src069[37] << 69) +
      (src069[38] << 69) +
      (src069[39] << 69) +
      (src069[40] << 69) +
      (src069[41] << 69) +
      (src069[42] << 69) +
      (src069[43] << 69) +
      (src069[44] << 69) +
      (src069[45] << 69) +
      (src069[46] << 69) +
      (src069[47] << 69) +
      (src069[48] << 69) +
      (src069[49] << 69) +
      (src069[50] << 69) +
      (src069[51] << 69) +
      (src069[52] << 69) +
      (src069[53] << 69) +
      (src069[54] << 69) +
      (src069[55] << 69) +
      (src069[56] << 69) +
      (src069[57] << 69) +
      (src069[58] << 69) +
      (src069[59] << 69) +
      (src069[60] << 69) +
      (src069[61] << 69) +
      (src069[62] << 69) +
      (src069[63] << 69) +
      (src069[64] << 69) +
      (src069[65] << 69) +
      (src069[66] << 69) +
      (src069[67] << 69) +
      (src069[68] << 69) +
      (src069[69] << 69) +
      (src069[70] << 69) +
      (src069[71] << 69) +
      (src069[72] << 69) +
      (src069[73] << 69) +
      (src069[74] << 69) +
      (src069[75] << 69) +
      (src069[76] << 69) +
      (src069[77] << 69) +
      (src069[78] << 69) +
      (src069[79] << 69) +
      (src069[80] << 69) +
      (src069[81] << 69) +
      (src069[82] << 69) +
      (src069[83] << 69) +
      (src069[84] << 69) +
      (src069[85] << 69) +
      (src069[86] << 69) +
      (src069[87] << 69) +
      (src069[88] << 69) +
      (src069[89] << 69) +
      (src069[90] << 69) +
      (src069[91] << 69) +
      (src069[92] << 69) +
      (src069[93] << 69) +
      (src069[94] << 69) +
      (src069[95] << 69) +
      (src069[96] << 69) +
      (src069[97] << 69) +
      (src069[98] << 69) +
      (src069[99] << 69) +
      (src069[100] << 69) +
      (src069[101] << 69) +
      (src069[102] << 69) +
      (src069[103] << 69) +
      (src069[104] << 69) +
      (src069[105] << 69) +
      (src069[106] << 69) +
      (src069[107] << 69) +
      (src069[108] << 69) +
      (src069[109] << 69) +
      (src069[110] << 69) +
      (src069[111] << 69) +
      (src069[112] << 69) +
      (src069[113] << 69) +
      (src069[114] << 69) +
      (src069[115] << 69) +
      (src069[116] << 69) +
      (src069[117] << 69) +
      (src069[118] << 69) +
      (src069[119] << 69) +
      (src069[120] << 69) +
      (src069[121] << 69) +
      (src069[122] << 69) +
      (src069[123] << 69) +
      (src069[124] << 69) +
      (src069[125] << 69) +
      (src069[126] << 69) +
      (src069[127] << 69) +
      (src070[0] << 70) +
      (src070[1] << 70) +
      (src070[2] << 70) +
      (src070[3] << 70) +
      (src070[4] << 70) +
      (src070[5] << 70) +
      (src070[6] << 70) +
      (src070[7] << 70) +
      (src070[8] << 70) +
      (src070[9] << 70) +
      (src070[10] << 70) +
      (src070[11] << 70) +
      (src070[12] << 70) +
      (src070[13] << 70) +
      (src070[14] << 70) +
      (src070[15] << 70) +
      (src070[16] << 70) +
      (src070[17] << 70) +
      (src070[18] << 70) +
      (src070[19] << 70) +
      (src070[20] << 70) +
      (src070[21] << 70) +
      (src070[22] << 70) +
      (src070[23] << 70) +
      (src070[24] << 70) +
      (src070[25] << 70) +
      (src070[26] << 70) +
      (src070[27] << 70) +
      (src070[28] << 70) +
      (src070[29] << 70) +
      (src070[30] << 70) +
      (src070[31] << 70) +
      (src070[32] << 70) +
      (src070[33] << 70) +
      (src070[34] << 70) +
      (src070[35] << 70) +
      (src070[36] << 70) +
      (src070[37] << 70) +
      (src070[38] << 70) +
      (src070[39] << 70) +
      (src070[40] << 70) +
      (src070[41] << 70) +
      (src070[42] << 70) +
      (src070[43] << 70) +
      (src070[44] << 70) +
      (src070[45] << 70) +
      (src070[46] << 70) +
      (src070[47] << 70) +
      (src070[48] << 70) +
      (src070[49] << 70) +
      (src070[50] << 70) +
      (src070[51] << 70) +
      (src070[52] << 70) +
      (src070[53] << 70) +
      (src070[54] << 70) +
      (src070[55] << 70) +
      (src070[56] << 70) +
      (src070[57] << 70) +
      (src070[58] << 70) +
      (src070[59] << 70) +
      (src070[60] << 70) +
      (src070[61] << 70) +
      (src070[62] << 70) +
      (src070[63] << 70) +
      (src070[64] << 70) +
      (src070[65] << 70) +
      (src070[66] << 70) +
      (src070[67] << 70) +
      (src070[68] << 70) +
      (src070[69] << 70) +
      (src070[70] << 70) +
      (src070[71] << 70) +
      (src070[72] << 70) +
      (src070[73] << 70) +
      (src070[74] << 70) +
      (src070[75] << 70) +
      (src070[76] << 70) +
      (src070[77] << 70) +
      (src070[78] << 70) +
      (src070[79] << 70) +
      (src070[80] << 70) +
      (src070[81] << 70) +
      (src070[82] << 70) +
      (src070[83] << 70) +
      (src070[84] << 70) +
      (src070[85] << 70) +
      (src070[86] << 70) +
      (src070[87] << 70) +
      (src070[88] << 70) +
      (src070[89] << 70) +
      (src070[90] << 70) +
      (src070[91] << 70) +
      (src070[92] << 70) +
      (src070[93] << 70) +
      (src070[94] << 70) +
      (src070[95] << 70) +
      (src070[96] << 70) +
      (src070[97] << 70) +
      (src070[98] << 70) +
      (src070[99] << 70) +
      (src070[100] << 70) +
      (src070[101] << 70) +
      (src070[102] << 70) +
      (src070[103] << 70) +
      (src070[104] << 70) +
      (src070[105] << 70) +
      (src070[106] << 70) +
      (src070[107] << 70) +
      (src070[108] << 70) +
      (src070[109] << 70) +
      (src070[110] << 70) +
      (src070[111] << 70) +
      (src070[112] << 70) +
      (src070[113] << 70) +
      (src070[114] << 70) +
      (src070[115] << 70) +
      (src070[116] << 70) +
      (src070[117] << 70) +
      (src070[118] << 70) +
      (src070[119] << 70) +
      (src070[120] << 70) +
      (src070[121] << 70) +
      (src070[122] << 70) +
      (src070[123] << 70) +
      (src070[124] << 70) +
      (src070[125] << 70) +
      (src070[126] << 70) +
      (src070[127] << 70) +
      (src071[0] << 71) +
      (src071[1] << 71) +
      (src071[2] << 71) +
      (src071[3] << 71) +
      (src071[4] << 71) +
      (src071[5] << 71) +
      (src071[6] << 71) +
      (src071[7] << 71) +
      (src071[8] << 71) +
      (src071[9] << 71) +
      (src071[10] << 71) +
      (src071[11] << 71) +
      (src071[12] << 71) +
      (src071[13] << 71) +
      (src071[14] << 71) +
      (src071[15] << 71) +
      (src071[16] << 71) +
      (src071[17] << 71) +
      (src071[18] << 71) +
      (src071[19] << 71) +
      (src071[20] << 71) +
      (src071[21] << 71) +
      (src071[22] << 71) +
      (src071[23] << 71) +
      (src071[24] << 71) +
      (src071[25] << 71) +
      (src071[26] << 71) +
      (src071[27] << 71) +
      (src071[28] << 71) +
      (src071[29] << 71) +
      (src071[30] << 71) +
      (src071[31] << 71) +
      (src071[32] << 71) +
      (src071[33] << 71) +
      (src071[34] << 71) +
      (src071[35] << 71) +
      (src071[36] << 71) +
      (src071[37] << 71) +
      (src071[38] << 71) +
      (src071[39] << 71) +
      (src071[40] << 71) +
      (src071[41] << 71) +
      (src071[42] << 71) +
      (src071[43] << 71) +
      (src071[44] << 71) +
      (src071[45] << 71) +
      (src071[46] << 71) +
      (src071[47] << 71) +
      (src071[48] << 71) +
      (src071[49] << 71) +
      (src071[50] << 71) +
      (src071[51] << 71) +
      (src071[52] << 71) +
      (src071[53] << 71) +
      (src071[54] << 71) +
      (src071[55] << 71) +
      (src071[56] << 71) +
      (src071[57] << 71) +
      (src071[58] << 71) +
      (src071[59] << 71) +
      (src071[60] << 71) +
      (src071[61] << 71) +
      (src071[62] << 71) +
      (src071[63] << 71) +
      (src071[64] << 71) +
      (src071[65] << 71) +
      (src071[66] << 71) +
      (src071[67] << 71) +
      (src071[68] << 71) +
      (src071[69] << 71) +
      (src071[70] << 71) +
      (src071[71] << 71) +
      (src071[72] << 71) +
      (src071[73] << 71) +
      (src071[74] << 71) +
      (src071[75] << 71) +
      (src071[76] << 71) +
      (src071[77] << 71) +
      (src071[78] << 71) +
      (src071[79] << 71) +
      (src071[80] << 71) +
      (src071[81] << 71) +
      (src071[82] << 71) +
      (src071[83] << 71) +
      (src071[84] << 71) +
      (src071[85] << 71) +
      (src071[86] << 71) +
      (src071[87] << 71) +
      (src071[88] << 71) +
      (src071[89] << 71) +
      (src071[90] << 71) +
      (src071[91] << 71) +
      (src071[92] << 71) +
      (src071[93] << 71) +
      (src071[94] << 71) +
      (src071[95] << 71) +
      (src071[96] << 71) +
      (src071[97] << 71) +
      (src071[98] << 71) +
      (src071[99] << 71) +
      (src071[100] << 71) +
      (src071[101] << 71) +
      (src071[102] << 71) +
      (src071[103] << 71) +
      (src071[104] << 71) +
      (src071[105] << 71) +
      (src071[106] << 71) +
      (src071[107] << 71) +
      (src071[108] << 71) +
      (src071[109] << 71) +
      (src071[110] << 71) +
      (src071[111] << 71) +
      (src071[112] << 71) +
      (src071[113] << 71) +
      (src071[114] << 71) +
      (src071[115] << 71) +
      (src071[116] << 71) +
      (src071[117] << 71) +
      (src071[118] << 71) +
      (src071[119] << 71) +
      (src071[120] << 71) +
      (src071[121] << 71) +
      (src071[122] << 71) +
      (src071[123] << 71) +
      (src071[124] << 71) +
      (src071[125] << 71) +
      (src071[126] << 71) +
      (src071[127] << 71) +
      (src072[0] << 72) +
      (src072[1] << 72) +
      (src072[2] << 72) +
      (src072[3] << 72) +
      (src072[4] << 72) +
      (src072[5] << 72) +
      (src072[6] << 72) +
      (src072[7] << 72) +
      (src072[8] << 72) +
      (src072[9] << 72) +
      (src072[10] << 72) +
      (src072[11] << 72) +
      (src072[12] << 72) +
      (src072[13] << 72) +
      (src072[14] << 72) +
      (src072[15] << 72) +
      (src072[16] << 72) +
      (src072[17] << 72) +
      (src072[18] << 72) +
      (src072[19] << 72) +
      (src072[20] << 72) +
      (src072[21] << 72) +
      (src072[22] << 72) +
      (src072[23] << 72) +
      (src072[24] << 72) +
      (src072[25] << 72) +
      (src072[26] << 72) +
      (src072[27] << 72) +
      (src072[28] << 72) +
      (src072[29] << 72) +
      (src072[30] << 72) +
      (src072[31] << 72) +
      (src072[32] << 72) +
      (src072[33] << 72) +
      (src072[34] << 72) +
      (src072[35] << 72) +
      (src072[36] << 72) +
      (src072[37] << 72) +
      (src072[38] << 72) +
      (src072[39] << 72) +
      (src072[40] << 72) +
      (src072[41] << 72) +
      (src072[42] << 72) +
      (src072[43] << 72) +
      (src072[44] << 72) +
      (src072[45] << 72) +
      (src072[46] << 72) +
      (src072[47] << 72) +
      (src072[48] << 72) +
      (src072[49] << 72) +
      (src072[50] << 72) +
      (src072[51] << 72) +
      (src072[52] << 72) +
      (src072[53] << 72) +
      (src072[54] << 72) +
      (src072[55] << 72) +
      (src072[56] << 72) +
      (src072[57] << 72) +
      (src072[58] << 72) +
      (src072[59] << 72) +
      (src072[60] << 72) +
      (src072[61] << 72) +
      (src072[62] << 72) +
      (src072[63] << 72) +
      (src072[64] << 72) +
      (src072[65] << 72) +
      (src072[66] << 72) +
      (src072[67] << 72) +
      (src072[68] << 72) +
      (src072[69] << 72) +
      (src072[70] << 72) +
      (src072[71] << 72) +
      (src072[72] << 72) +
      (src072[73] << 72) +
      (src072[74] << 72) +
      (src072[75] << 72) +
      (src072[76] << 72) +
      (src072[77] << 72) +
      (src072[78] << 72) +
      (src072[79] << 72) +
      (src072[80] << 72) +
      (src072[81] << 72) +
      (src072[82] << 72) +
      (src072[83] << 72) +
      (src072[84] << 72) +
      (src072[85] << 72) +
      (src072[86] << 72) +
      (src072[87] << 72) +
      (src072[88] << 72) +
      (src072[89] << 72) +
      (src072[90] << 72) +
      (src072[91] << 72) +
      (src072[92] << 72) +
      (src072[93] << 72) +
      (src072[94] << 72) +
      (src072[95] << 72) +
      (src072[96] << 72) +
      (src072[97] << 72) +
      (src072[98] << 72) +
      (src072[99] << 72) +
      (src072[100] << 72) +
      (src072[101] << 72) +
      (src072[102] << 72) +
      (src072[103] << 72) +
      (src072[104] << 72) +
      (src072[105] << 72) +
      (src072[106] << 72) +
      (src072[107] << 72) +
      (src072[108] << 72) +
      (src072[109] << 72) +
      (src072[110] << 72) +
      (src072[111] << 72) +
      (src072[112] << 72) +
      (src072[113] << 72) +
      (src072[114] << 72) +
      (src072[115] << 72) +
      (src072[116] << 72) +
      (src072[117] << 72) +
      (src072[118] << 72) +
      (src072[119] << 72) +
      (src072[120] << 72) +
      (src072[121] << 72) +
      (src072[122] << 72) +
      (src072[123] << 72) +
      (src072[124] << 72) +
      (src072[125] << 72) +
      (src072[126] << 72) +
      (src072[127] << 72) +
      (src073[0] << 73) +
      (src073[1] << 73) +
      (src073[2] << 73) +
      (src073[3] << 73) +
      (src073[4] << 73) +
      (src073[5] << 73) +
      (src073[6] << 73) +
      (src073[7] << 73) +
      (src073[8] << 73) +
      (src073[9] << 73) +
      (src073[10] << 73) +
      (src073[11] << 73) +
      (src073[12] << 73) +
      (src073[13] << 73) +
      (src073[14] << 73) +
      (src073[15] << 73) +
      (src073[16] << 73) +
      (src073[17] << 73) +
      (src073[18] << 73) +
      (src073[19] << 73) +
      (src073[20] << 73) +
      (src073[21] << 73) +
      (src073[22] << 73) +
      (src073[23] << 73) +
      (src073[24] << 73) +
      (src073[25] << 73) +
      (src073[26] << 73) +
      (src073[27] << 73) +
      (src073[28] << 73) +
      (src073[29] << 73) +
      (src073[30] << 73) +
      (src073[31] << 73) +
      (src073[32] << 73) +
      (src073[33] << 73) +
      (src073[34] << 73) +
      (src073[35] << 73) +
      (src073[36] << 73) +
      (src073[37] << 73) +
      (src073[38] << 73) +
      (src073[39] << 73) +
      (src073[40] << 73) +
      (src073[41] << 73) +
      (src073[42] << 73) +
      (src073[43] << 73) +
      (src073[44] << 73) +
      (src073[45] << 73) +
      (src073[46] << 73) +
      (src073[47] << 73) +
      (src073[48] << 73) +
      (src073[49] << 73) +
      (src073[50] << 73) +
      (src073[51] << 73) +
      (src073[52] << 73) +
      (src073[53] << 73) +
      (src073[54] << 73) +
      (src073[55] << 73) +
      (src073[56] << 73) +
      (src073[57] << 73) +
      (src073[58] << 73) +
      (src073[59] << 73) +
      (src073[60] << 73) +
      (src073[61] << 73) +
      (src073[62] << 73) +
      (src073[63] << 73) +
      (src073[64] << 73) +
      (src073[65] << 73) +
      (src073[66] << 73) +
      (src073[67] << 73) +
      (src073[68] << 73) +
      (src073[69] << 73) +
      (src073[70] << 73) +
      (src073[71] << 73) +
      (src073[72] << 73) +
      (src073[73] << 73) +
      (src073[74] << 73) +
      (src073[75] << 73) +
      (src073[76] << 73) +
      (src073[77] << 73) +
      (src073[78] << 73) +
      (src073[79] << 73) +
      (src073[80] << 73) +
      (src073[81] << 73) +
      (src073[82] << 73) +
      (src073[83] << 73) +
      (src073[84] << 73) +
      (src073[85] << 73) +
      (src073[86] << 73) +
      (src073[87] << 73) +
      (src073[88] << 73) +
      (src073[89] << 73) +
      (src073[90] << 73) +
      (src073[91] << 73) +
      (src073[92] << 73) +
      (src073[93] << 73) +
      (src073[94] << 73) +
      (src073[95] << 73) +
      (src073[96] << 73) +
      (src073[97] << 73) +
      (src073[98] << 73) +
      (src073[99] << 73) +
      (src073[100] << 73) +
      (src073[101] << 73) +
      (src073[102] << 73) +
      (src073[103] << 73) +
      (src073[104] << 73) +
      (src073[105] << 73) +
      (src073[106] << 73) +
      (src073[107] << 73) +
      (src073[108] << 73) +
      (src073[109] << 73) +
      (src073[110] << 73) +
      (src073[111] << 73) +
      (src073[112] << 73) +
      (src073[113] << 73) +
      (src073[114] << 73) +
      (src073[115] << 73) +
      (src073[116] << 73) +
      (src073[117] << 73) +
      (src073[118] << 73) +
      (src073[119] << 73) +
      (src073[120] << 73) +
      (src073[121] << 73) +
      (src073[122] << 73) +
      (src073[123] << 73) +
      (src073[124] << 73) +
      (src073[125] << 73) +
      (src073[126] << 73) +
      (src073[127] << 73) +
      (src074[0] << 74) +
      (src074[1] << 74) +
      (src074[2] << 74) +
      (src074[3] << 74) +
      (src074[4] << 74) +
      (src074[5] << 74) +
      (src074[6] << 74) +
      (src074[7] << 74) +
      (src074[8] << 74) +
      (src074[9] << 74) +
      (src074[10] << 74) +
      (src074[11] << 74) +
      (src074[12] << 74) +
      (src074[13] << 74) +
      (src074[14] << 74) +
      (src074[15] << 74) +
      (src074[16] << 74) +
      (src074[17] << 74) +
      (src074[18] << 74) +
      (src074[19] << 74) +
      (src074[20] << 74) +
      (src074[21] << 74) +
      (src074[22] << 74) +
      (src074[23] << 74) +
      (src074[24] << 74) +
      (src074[25] << 74) +
      (src074[26] << 74) +
      (src074[27] << 74) +
      (src074[28] << 74) +
      (src074[29] << 74) +
      (src074[30] << 74) +
      (src074[31] << 74) +
      (src074[32] << 74) +
      (src074[33] << 74) +
      (src074[34] << 74) +
      (src074[35] << 74) +
      (src074[36] << 74) +
      (src074[37] << 74) +
      (src074[38] << 74) +
      (src074[39] << 74) +
      (src074[40] << 74) +
      (src074[41] << 74) +
      (src074[42] << 74) +
      (src074[43] << 74) +
      (src074[44] << 74) +
      (src074[45] << 74) +
      (src074[46] << 74) +
      (src074[47] << 74) +
      (src074[48] << 74) +
      (src074[49] << 74) +
      (src074[50] << 74) +
      (src074[51] << 74) +
      (src074[52] << 74) +
      (src074[53] << 74) +
      (src074[54] << 74) +
      (src074[55] << 74) +
      (src074[56] << 74) +
      (src074[57] << 74) +
      (src074[58] << 74) +
      (src074[59] << 74) +
      (src074[60] << 74) +
      (src074[61] << 74) +
      (src074[62] << 74) +
      (src074[63] << 74) +
      (src074[64] << 74) +
      (src074[65] << 74) +
      (src074[66] << 74) +
      (src074[67] << 74) +
      (src074[68] << 74) +
      (src074[69] << 74) +
      (src074[70] << 74) +
      (src074[71] << 74) +
      (src074[72] << 74) +
      (src074[73] << 74) +
      (src074[74] << 74) +
      (src074[75] << 74) +
      (src074[76] << 74) +
      (src074[77] << 74) +
      (src074[78] << 74) +
      (src074[79] << 74) +
      (src074[80] << 74) +
      (src074[81] << 74) +
      (src074[82] << 74) +
      (src074[83] << 74) +
      (src074[84] << 74) +
      (src074[85] << 74) +
      (src074[86] << 74) +
      (src074[87] << 74) +
      (src074[88] << 74) +
      (src074[89] << 74) +
      (src074[90] << 74) +
      (src074[91] << 74) +
      (src074[92] << 74) +
      (src074[93] << 74) +
      (src074[94] << 74) +
      (src074[95] << 74) +
      (src074[96] << 74) +
      (src074[97] << 74) +
      (src074[98] << 74) +
      (src074[99] << 74) +
      (src074[100] << 74) +
      (src074[101] << 74) +
      (src074[102] << 74) +
      (src074[103] << 74) +
      (src074[104] << 74) +
      (src074[105] << 74) +
      (src074[106] << 74) +
      (src074[107] << 74) +
      (src074[108] << 74) +
      (src074[109] << 74) +
      (src074[110] << 74) +
      (src074[111] << 74) +
      (src074[112] << 74) +
      (src074[113] << 74) +
      (src074[114] << 74) +
      (src074[115] << 74) +
      (src074[116] << 74) +
      (src074[117] << 74) +
      (src074[118] << 74) +
      (src074[119] << 74) +
      (src074[120] << 74) +
      (src074[121] << 74) +
      (src074[122] << 74) +
      (src074[123] << 74) +
      (src074[124] << 74) +
      (src074[125] << 74) +
      (src074[126] << 74) +
      (src074[127] << 74) +
      (src075[0] << 75) +
      (src075[1] << 75) +
      (src075[2] << 75) +
      (src075[3] << 75) +
      (src075[4] << 75) +
      (src075[5] << 75) +
      (src075[6] << 75) +
      (src075[7] << 75) +
      (src075[8] << 75) +
      (src075[9] << 75) +
      (src075[10] << 75) +
      (src075[11] << 75) +
      (src075[12] << 75) +
      (src075[13] << 75) +
      (src075[14] << 75) +
      (src075[15] << 75) +
      (src075[16] << 75) +
      (src075[17] << 75) +
      (src075[18] << 75) +
      (src075[19] << 75) +
      (src075[20] << 75) +
      (src075[21] << 75) +
      (src075[22] << 75) +
      (src075[23] << 75) +
      (src075[24] << 75) +
      (src075[25] << 75) +
      (src075[26] << 75) +
      (src075[27] << 75) +
      (src075[28] << 75) +
      (src075[29] << 75) +
      (src075[30] << 75) +
      (src075[31] << 75) +
      (src075[32] << 75) +
      (src075[33] << 75) +
      (src075[34] << 75) +
      (src075[35] << 75) +
      (src075[36] << 75) +
      (src075[37] << 75) +
      (src075[38] << 75) +
      (src075[39] << 75) +
      (src075[40] << 75) +
      (src075[41] << 75) +
      (src075[42] << 75) +
      (src075[43] << 75) +
      (src075[44] << 75) +
      (src075[45] << 75) +
      (src075[46] << 75) +
      (src075[47] << 75) +
      (src075[48] << 75) +
      (src075[49] << 75) +
      (src075[50] << 75) +
      (src075[51] << 75) +
      (src075[52] << 75) +
      (src075[53] << 75) +
      (src075[54] << 75) +
      (src075[55] << 75) +
      (src075[56] << 75) +
      (src075[57] << 75) +
      (src075[58] << 75) +
      (src075[59] << 75) +
      (src075[60] << 75) +
      (src075[61] << 75) +
      (src075[62] << 75) +
      (src075[63] << 75) +
      (src075[64] << 75) +
      (src075[65] << 75) +
      (src075[66] << 75) +
      (src075[67] << 75) +
      (src075[68] << 75) +
      (src075[69] << 75) +
      (src075[70] << 75) +
      (src075[71] << 75) +
      (src075[72] << 75) +
      (src075[73] << 75) +
      (src075[74] << 75) +
      (src075[75] << 75) +
      (src075[76] << 75) +
      (src075[77] << 75) +
      (src075[78] << 75) +
      (src075[79] << 75) +
      (src075[80] << 75) +
      (src075[81] << 75) +
      (src075[82] << 75) +
      (src075[83] << 75) +
      (src075[84] << 75) +
      (src075[85] << 75) +
      (src075[86] << 75) +
      (src075[87] << 75) +
      (src075[88] << 75) +
      (src075[89] << 75) +
      (src075[90] << 75) +
      (src075[91] << 75) +
      (src075[92] << 75) +
      (src075[93] << 75) +
      (src075[94] << 75) +
      (src075[95] << 75) +
      (src075[96] << 75) +
      (src075[97] << 75) +
      (src075[98] << 75) +
      (src075[99] << 75) +
      (src075[100] << 75) +
      (src075[101] << 75) +
      (src075[102] << 75) +
      (src075[103] << 75) +
      (src075[104] << 75) +
      (src075[105] << 75) +
      (src075[106] << 75) +
      (src075[107] << 75) +
      (src075[108] << 75) +
      (src075[109] << 75) +
      (src075[110] << 75) +
      (src075[111] << 75) +
      (src075[112] << 75) +
      (src075[113] << 75) +
      (src075[114] << 75) +
      (src075[115] << 75) +
      (src075[116] << 75) +
      (src075[117] << 75) +
      (src075[118] << 75) +
      (src075[119] << 75) +
      (src075[120] << 75) +
      (src075[121] << 75) +
      (src075[122] << 75) +
      (src075[123] << 75) +
      (src075[124] << 75) +
      (src075[125] << 75) +
      (src075[126] << 75) +
      (src075[127] << 75) +
      (src076[0] << 76) +
      (src076[1] << 76) +
      (src076[2] << 76) +
      (src076[3] << 76) +
      (src076[4] << 76) +
      (src076[5] << 76) +
      (src076[6] << 76) +
      (src076[7] << 76) +
      (src076[8] << 76) +
      (src076[9] << 76) +
      (src076[10] << 76) +
      (src076[11] << 76) +
      (src076[12] << 76) +
      (src076[13] << 76) +
      (src076[14] << 76) +
      (src076[15] << 76) +
      (src076[16] << 76) +
      (src076[17] << 76) +
      (src076[18] << 76) +
      (src076[19] << 76) +
      (src076[20] << 76) +
      (src076[21] << 76) +
      (src076[22] << 76) +
      (src076[23] << 76) +
      (src076[24] << 76) +
      (src076[25] << 76) +
      (src076[26] << 76) +
      (src076[27] << 76) +
      (src076[28] << 76) +
      (src076[29] << 76) +
      (src076[30] << 76) +
      (src076[31] << 76) +
      (src076[32] << 76) +
      (src076[33] << 76) +
      (src076[34] << 76) +
      (src076[35] << 76) +
      (src076[36] << 76) +
      (src076[37] << 76) +
      (src076[38] << 76) +
      (src076[39] << 76) +
      (src076[40] << 76) +
      (src076[41] << 76) +
      (src076[42] << 76) +
      (src076[43] << 76) +
      (src076[44] << 76) +
      (src076[45] << 76) +
      (src076[46] << 76) +
      (src076[47] << 76) +
      (src076[48] << 76) +
      (src076[49] << 76) +
      (src076[50] << 76) +
      (src076[51] << 76) +
      (src076[52] << 76) +
      (src076[53] << 76) +
      (src076[54] << 76) +
      (src076[55] << 76) +
      (src076[56] << 76) +
      (src076[57] << 76) +
      (src076[58] << 76) +
      (src076[59] << 76) +
      (src076[60] << 76) +
      (src076[61] << 76) +
      (src076[62] << 76) +
      (src076[63] << 76) +
      (src076[64] << 76) +
      (src076[65] << 76) +
      (src076[66] << 76) +
      (src076[67] << 76) +
      (src076[68] << 76) +
      (src076[69] << 76) +
      (src076[70] << 76) +
      (src076[71] << 76) +
      (src076[72] << 76) +
      (src076[73] << 76) +
      (src076[74] << 76) +
      (src076[75] << 76) +
      (src076[76] << 76) +
      (src076[77] << 76) +
      (src076[78] << 76) +
      (src076[79] << 76) +
      (src076[80] << 76) +
      (src076[81] << 76) +
      (src076[82] << 76) +
      (src076[83] << 76) +
      (src076[84] << 76) +
      (src076[85] << 76) +
      (src076[86] << 76) +
      (src076[87] << 76) +
      (src076[88] << 76) +
      (src076[89] << 76) +
      (src076[90] << 76) +
      (src076[91] << 76) +
      (src076[92] << 76) +
      (src076[93] << 76) +
      (src076[94] << 76) +
      (src076[95] << 76) +
      (src076[96] << 76) +
      (src076[97] << 76) +
      (src076[98] << 76) +
      (src076[99] << 76) +
      (src076[100] << 76) +
      (src076[101] << 76) +
      (src076[102] << 76) +
      (src076[103] << 76) +
      (src076[104] << 76) +
      (src076[105] << 76) +
      (src076[106] << 76) +
      (src076[107] << 76) +
      (src076[108] << 76) +
      (src076[109] << 76) +
      (src076[110] << 76) +
      (src076[111] << 76) +
      (src076[112] << 76) +
      (src076[113] << 76) +
      (src076[114] << 76) +
      (src076[115] << 76) +
      (src076[116] << 76) +
      (src076[117] << 76) +
      (src076[118] << 76) +
      (src076[119] << 76) +
      (src076[120] << 76) +
      (src076[121] << 76) +
      (src076[122] << 76) +
      (src076[123] << 76) +
      (src076[124] << 76) +
      (src076[125] << 76) +
      (src076[126] << 76) +
      (src076[127] << 76) +
      (src077[0] << 77) +
      (src077[1] << 77) +
      (src077[2] << 77) +
      (src077[3] << 77) +
      (src077[4] << 77) +
      (src077[5] << 77) +
      (src077[6] << 77) +
      (src077[7] << 77) +
      (src077[8] << 77) +
      (src077[9] << 77) +
      (src077[10] << 77) +
      (src077[11] << 77) +
      (src077[12] << 77) +
      (src077[13] << 77) +
      (src077[14] << 77) +
      (src077[15] << 77) +
      (src077[16] << 77) +
      (src077[17] << 77) +
      (src077[18] << 77) +
      (src077[19] << 77) +
      (src077[20] << 77) +
      (src077[21] << 77) +
      (src077[22] << 77) +
      (src077[23] << 77) +
      (src077[24] << 77) +
      (src077[25] << 77) +
      (src077[26] << 77) +
      (src077[27] << 77) +
      (src077[28] << 77) +
      (src077[29] << 77) +
      (src077[30] << 77) +
      (src077[31] << 77) +
      (src077[32] << 77) +
      (src077[33] << 77) +
      (src077[34] << 77) +
      (src077[35] << 77) +
      (src077[36] << 77) +
      (src077[37] << 77) +
      (src077[38] << 77) +
      (src077[39] << 77) +
      (src077[40] << 77) +
      (src077[41] << 77) +
      (src077[42] << 77) +
      (src077[43] << 77) +
      (src077[44] << 77) +
      (src077[45] << 77) +
      (src077[46] << 77) +
      (src077[47] << 77) +
      (src077[48] << 77) +
      (src077[49] << 77) +
      (src077[50] << 77) +
      (src077[51] << 77) +
      (src077[52] << 77) +
      (src077[53] << 77) +
      (src077[54] << 77) +
      (src077[55] << 77) +
      (src077[56] << 77) +
      (src077[57] << 77) +
      (src077[58] << 77) +
      (src077[59] << 77) +
      (src077[60] << 77) +
      (src077[61] << 77) +
      (src077[62] << 77) +
      (src077[63] << 77) +
      (src077[64] << 77) +
      (src077[65] << 77) +
      (src077[66] << 77) +
      (src077[67] << 77) +
      (src077[68] << 77) +
      (src077[69] << 77) +
      (src077[70] << 77) +
      (src077[71] << 77) +
      (src077[72] << 77) +
      (src077[73] << 77) +
      (src077[74] << 77) +
      (src077[75] << 77) +
      (src077[76] << 77) +
      (src077[77] << 77) +
      (src077[78] << 77) +
      (src077[79] << 77) +
      (src077[80] << 77) +
      (src077[81] << 77) +
      (src077[82] << 77) +
      (src077[83] << 77) +
      (src077[84] << 77) +
      (src077[85] << 77) +
      (src077[86] << 77) +
      (src077[87] << 77) +
      (src077[88] << 77) +
      (src077[89] << 77) +
      (src077[90] << 77) +
      (src077[91] << 77) +
      (src077[92] << 77) +
      (src077[93] << 77) +
      (src077[94] << 77) +
      (src077[95] << 77) +
      (src077[96] << 77) +
      (src077[97] << 77) +
      (src077[98] << 77) +
      (src077[99] << 77) +
      (src077[100] << 77) +
      (src077[101] << 77) +
      (src077[102] << 77) +
      (src077[103] << 77) +
      (src077[104] << 77) +
      (src077[105] << 77) +
      (src077[106] << 77) +
      (src077[107] << 77) +
      (src077[108] << 77) +
      (src077[109] << 77) +
      (src077[110] << 77) +
      (src077[111] << 77) +
      (src077[112] << 77) +
      (src077[113] << 77) +
      (src077[114] << 77) +
      (src077[115] << 77) +
      (src077[116] << 77) +
      (src077[117] << 77) +
      (src077[118] << 77) +
      (src077[119] << 77) +
      (src077[120] << 77) +
      (src077[121] << 77) +
      (src077[122] << 77) +
      (src077[123] << 77) +
      (src077[124] << 77) +
      (src077[125] << 77) +
      (src077[126] << 77) +
      (src077[127] << 77) +
      (src078[0] << 78) +
      (src078[1] << 78) +
      (src078[2] << 78) +
      (src078[3] << 78) +
      (src078[4] << 78) +
      (src078[5] << 78) +
      (src078[6] << 78) +
      (src078[7] << 78) +
      (src078[8] << 78) +
      (src078[9] << 78) +
      (src078[10] << 78) +
      (src078[11] << 78) +
      (src078[12] << 78) +
      (src078[13] << 78) +
      (src078[14] << 78) +
      (src078[15] << 78) +
      (src078[16] << 78) +
      (src078[17] << 78) +
      (src078[18] << 78) +
      (src078[19] << 78) +
      (src078[20] << 78) +
      (src078[21] << 78) +
      (src078[22] << 78) +
      (src078[23] << 78) +
      (src078[24] << 78) +
      (src078[25] << 78) +
      (src078[26] << 78) +
      (src078[27] << 78) +
      (src078[28] << 78) +
      (src078[29] << 78) +
      (src078[30] << 78) +
      (src078[31] << 78) +
      (src078[32] << 78) +
      (src078[33] << 78) +
      (src078[34] << 78) +
      (src078[35] << 78) +
      (src078[36] << 78) +
      (src078[37] << 78) +
      (src078[38] << 78) +
      (src078[39] << 78) +
      (src078[40] << 78) +
      (src078[41] << 78) +
      (src078[42] << 78) +
      (src078[43] << 78) +
      (src078[44] << 78) +
      (src078[45] << 78) +
      (src078[46] << 78) +
      (src078[47] << 78) +
      (src078[48] << 78) +
      (src078[49] << 78) +
      (src078[50] << 78) +
      (src078[51] << 78) +
      (src078[52] << 78) +
      (src078[53] << 78) +
      (src078[54] << 78) +
      (src078[55] << 78) +
      (src078[56] << 78) +
      (src078[57] << 78) +
      (src078[58] << 78) +
      (src078[59] << 78) +
      (src078[60] << 78) +
      (src078[61] << 78) +
      (src078[62] << 78) +
      (src078[63] << 78) +
      (src078[64] << 78) +
      (src078[65] << 78) +
      (src078[66] << 78) +
      (src078[67] << 78) +
      (src078[68] << 78) +
      (src078[69] << 78) +
      (src078[70] << 78) +
      (src078[71] << 78) +
      (src078[72] << 78) +
      (src078[73] << 78) +
      (src078[74] << 78) +
      (src078[75] << 78) +
      (src078[76] << 78) +
      (src078[77] << 78) +
      (src078[78] << 78) +
      (src078[79] << 78) +
      (src078[80] << 78) +
      (src078[81] << 78) +
      (src078[82] << 78) +
      (src078[83] << 78) +
      (src078[84] << 78) +
      (src078[85] << 78) +
      (src078[86] << 78) +
      (src078[87] << 78) +
      (src078[88] << 78) +
      (src078[89] << 78) +
      (src078[90] << 78) +
      (src078[91] << 78) +
      (src078[92] << 78) +
      (src078[93] << 78) +
      (src078[94] << 78) +
      (src078[95] << 78) +
      (src078[96] << 78) +
      (src078[97] << 78) +
      (src078[98] << 78) +
      (src078[99] << 78) +
      (src078[100] << 78) +
      (src078[101] << 78) +
      (src078[102] << 78) +
      (src078[103] << 78) +
      (src078[104] << 78) +
      (src078[105] << 78) +
      (src078[106] << 78) +
      (src078[107] << 78) +
      (src078[108] << 78) +
      (src078[109] << 78) +
      (src078[110] << 78) +
      (src078[111] << 78) +
      (src078[112] << 78) +
      (src078[113] << 78) +
      (src078[114] << 78) +
      (src078[115] << 78) +
      (src078[116] << 78) +
      (src078[117] << 78) +
      (src078[118] << 78) +
      (src078[119] << 78) +
      (src078[120] << 78) +
      (src078[121] << 78) +
      (src078[122] << 78) +
      (src078[123] << 78) +
      (src078[124] << 78) +
      (src078[125] << 78) +
      (src078[126] << 78) +
      (src078[127] << 78) +
      (src079[0] << 79) +
      (src079[1] << 79) +
      (src079[2] << 79) +
      (src079[3] << 79) +
      (src079[4] << 79) +
      (src079[5] << 79) +
      (src079[6] << 79) +
      (src079[7] << 79) +
      (src079[8] << 79) +
      (src079[9] << 79) +
      (src079[10] << 79) +
      (src079[11] << 79) +
      (src079[12] << 79) +
      (src079[13] << 79) +
      (src079[14] << 79) +
      (src079[15] << 79) +
      (src079[16] << 79) +
      (src079[17] << 79) +
      (src079[18] << 79) +
      (src079[19] << 79) +
      (src079[20] << 79) +
      (src079[21] << 79) +
      (src079[22] << 79) +
      (src079[23] << 79) +
      (src079[24] << 79) +
      (src079[25] << 79) +
      (src079[26] << 79) +
      (src079[27] << 79) +
      (src079[28] << 79) +
      (src079[29] << 79) +
      (src079[30] << 79) +
      (src079[31] << 79) +
      (src079[32] << 79) +
      (src079[33] << 79) +
      (src079[34] << 79) +
      (src079[35] << 79) +
      (src079[36] << 79) +
      (src079[37] << 79) +
      (src079[38] << 79) +
      (src079[39] << 79) +
      (src079[40] << 79) +
      (src079[41] << 79) +
      (src079[42] << 79) +
      (src079[43] << 79) +
      (src079[44] << 79) +
      (src079[45] << 79) +
      (src079[46] << 79) +
      (src079[47] << 79) +
      (src079[48] << 79) +
      (src079[49] << 79) +
      (src079[50] << 79) +
      (src079[51] << 79) +
      (src079[52] << 79) +
      (src079[53] << 79) +
      (src079[54] << 79) +
      (src079[55] << 79) +
      (src079[56] << 79) +
      (src079[57] << 79) +
      (src079[58] << 79) +
      (src079[59] << 79) +
      (src079[60] << 79) +
      (src079[61] << 79) +
      (src079[62] << 79) +
      (src079[63] << 79) +
      (src079[64] << 79) +
      (src079[65] << 79) +
      (src079[66] << 79) +
      (src079[67] << 79) +
      (src079[68] << 79) +
      (src079[69] << 79) +
      (src079[70] << 79) +
      (src079[71] << 79) +
      (src079[72] << 79) +
      (src079[73] << 79) +
      (src079[74] << 79) +
      (src079[75] << 79) +
      (src079[76] << 79) +
      (src079[77] << 79) +
      (src079[78] << 79) +
      (src079[79] << 79) +
      (src079[80] << 79) +
      (src079[81] << 79) +
      (src079[82] << 79) +
      (src079[83] << 79) +
      (src079[84] << 79) +
      (src079[85] << 79) +
      (src079[86] << 79) +
      (src079[87] << 79) +
      (src079[88] << 79) +
      (src079[89] << 79) +
      (src079[90] << 79) +
      (src079[91] << 79) +
      (src079[92] << 79) +
      (src079[93] << 79) +
      (src079[94] << 79) +
      (src079[95] << 79) +
      (src079[96] << 79) +
      (src079[97] << 79) +
      (src079[98] << 79) +
      (src079[99] << 79) +
      (src079[100] << 79) +
      (src079[101] << 79) +
      (src079[102] << 79) +
      (src079[103] << 79) +
      (src079[104] << 79) +
      (src079[105] << 79) +
      (src079[106] << 79) +
      (src079[107] << 79) +
      (src079[108] << 79) +
      (src079[109] << 79) +
      (src079[110] << 79) +
      (src079[111] << 79) +
      (src079[112] << 79) +
      (src079[113] << 79) +
      (src079[114] << 79) +
      (src079[115] << 79) +
      (src079[116] << 79) +
      (src079[117] << 79) +
      (src079[118] << 79) +
      (src079[119] << 79) +
      (src079[120] << 79) +
      (src079[121] << 79) +
      (src079[122] << 79) +
      (src079[123] << 79) +
      (src079[124] << 79) +
      (src079[125] << 79) +
      (src079[126] << 79) +
      (src079[127] << 79) +
      (src080[0] << 80) +
      (src080[1] << 80) +
      (src080[2] << 80) +
      (src080[3] << 80) +
      (src080[4] << 80) +
      (src080[5] << 80) +
      (src080[6] << 80) +
      (src080[7] << 80) +
      (src080[8] << 80) +
      (src080[9] << 80) +
      (src080[10] << 80) +
      (src080[11] << 80) +
      (src080[12] << 80) +
      (src080[13] << 80) +
      (src080[14] << 80) +
      (src080[15] << 80) +
      (src080[16] << 80) +
      (src080[17] << 80) +
      (src080[18] << 80) +
      (src080[19] << 80) +
      (src080[20] << 80) +
      (src080[21] << 80) +
      (src080[22] << 80) +
      (src080[23] << 80) +
      (src080[24] << 80) +
      (src080[25] << 80) +
      (src080[26] << 80) +
      (src080[27] << 80) +
      (src080[28] << 80) +
      (src080[29] << 80) +
      (src080[30] << 80) +
      (src080[31] << 80) +
      (src080[32] << 80) +
      (src080[33] << 80) +
      (src080[34] << 80) +
      (src080[35] << 80) +
      (src080[36] << 80) +
      (src080[37] << 80) +
      (src080[38] << 80) +
      (src080[39] << 80) +
      (src080[40] << 80) +
      (src080[41] << 80) +
      (src080[42] << 80) +
      (src080[43] << 80) +
      (src080[44] << 80) +
      (src080[45] << 80) +
      (src080[46] << 80) +
      (src080[47] << 80) +
      (src080[48] << 80) +
      (src080[49] << 80) +
      (src080[50] << 80) +
      (src080[51] << 80) +
      (src080[52] << 80) +
      (src080[53] << 80) +
      (src080[54] << 80) +
      (src080[55] << 80) +
      (src080[56] << 80) +
      (src080[57] << 80) +
      (src080[58] << 80) +
      (src080[59] << 80) +
      (src080[60] << 80) +
      (src080[61] << 80) +
      (src080[62] << 80) +
      (src080[63] << 80) +
      (src080[64] << 80) +
      (src080[65] << 80) +
      (src080[66] << 80) +
      (src080[67] << 80) +
      (src080[68] << 80) +
      (src080[69] << 80) +
      (src080[70] << 80) +
      (src080[71] << 80) +
      (src080[72] << 80) +
      (src080[73] << 80) +
      (src080[74] << 80) +
      (src080[75] << 80) +
      (src080[76] << 80) +
      (src080[77] << 80) +
      (src080[78] << 80) +
      (src080[79] << 80) +
      (src080[80] << 80) +
      (src080[81] << 80) +
      (src080[82] << 80) +
      (src080[83] << 80) +
      (src080[84] << 80) +
      (src080[85] << 80) +
      (src080[86] << 80) +
      (src080[87] << 80) +
      (src080[88] << 80) +
      (src080[89] << 80) +
      (src080[90] << 80) +
      (src080[91] << 80) +
      (src080[92] << 80) +
      (src080[93] << 80) +
      (src080[94] << 80) +
      (src080[95] << 80) +
      (src080[96] << 80) +
      (src080[97] << 80) +
      (src080[98] << 80) +
      (src080[99] << 80) +
      (src080[100] << 80) +
      (src080[101] << 80) +
      (src080[102] << 80) +
      (src080[103] << 80) +
      (src080[104] << 80) +
      (src080[105] << 80) +
      (src080[106] << 80) +
      (src080[107] << 80) +
      (src080[108] << 80) +
      (src080[109] << 80) +
      (src080[110] << 80) +
      (src080[111] << 80) +
      (src080[112] << 80) +
      (src080[113] << 80) +
      (src080[114] << 80) +
      (src080[115] << 80) +
      (src080[116] << 80) +
      (src080[117] << 80) +
      (src080[118] << 80) +
      (src080[119] << 80) +
      (src080[120] << 80) +
      (src080[121] << 80) +
      (src080[122] << 80) +
      (src080[123] << 80) +
      (src080[124] << 80) +
      (src080[125] << 80) +
      (src080[126] << 80) +
      (src080[127] << 80) +
      (src081[0] << 81) +
      (src081[1] << 81) +
      (src081[2] << 81) +
      (src081[3] << 81) +
      (src081[4] << 81) +
      (src081[5] << 81) +
      (src081[6] << 81) +
      (src081[7] << 81) +
      (src081[8] << 81) +
      (src081[9] << 81) +
      (src081[10] << 81) +
      (src081[11] << 81) +
      (src081[12] << 81) +
      (src081[13] << 81) +
      (src081[14] << 81) +
      (src081[15] << 81) +
      (src081[16] << 81) +
      (src081[17] << 81) +
      (src081[18] << 81) +
      (src081[19] << 81) +
      (src081[20] << 81) +
      (src081[21] << 81) +
      (src081[22] << 81) +
      (src081[23] << 81) +
      (src081[24] << 81) +
      (src081[25] << 81) +
      (src081[26] << 81) +
      (src081[27] << 81) +
      (src081[28] << 81) +
      (src081[29] << 81) +
      (src081[30] << 81) +
      (src081[31] << 81) +
      (src081[32] << 81) +
      (src081[33] << 81) +
      (src081[34] << 81) +
      (src081[35] << 81) +
      (src081[36] << 81) +
      (src081[37] << 81) +
      (src081[38] << 81) +
      (src081[39] << 81) +
      (src081[40] << 81) +
      (src081[41] << 81) +
      (src081[42] << 81) +
      (src081[43] << 81) +
      (src081[44] << 81) +
      (src081[45] << 81) +
      (src081[46] << 81) +
      (src081[47] << 81) +
      (src081[48] << 81) +
      (src081[49] << 81) +
      (src081[50] << 81) +
      (src081[51] << 81) +
      (src081[52] << 81) +
      (src081[53] << 81) +
      (src081[54] << 81) +
      (src081[55] << 81) +
      (src081[56] << 81) +
      (src081[57] << 81) +
      (src081[58] << 81) +
      (src081[59] << 81) +
      (src081[60] << 81) +
      (src081[61] << 81) +
      (src081[62] << 81) +
      (src081[63] << 81) +
      (src081[64] << 81) +
      (src081[65] << 81) +
      (src081[66] << 81) +
      (src081[67] << 81) +
      (src081[68] << 81) +
      (src081[69] << 81) +
      (src081[70] << 81) +
      (src081[71] << 81) +
      (src081[72] << 81) +
      (src081[73] << 81) +
      (src081[74] << 81) +
      (src081[75] << 81) +
      (src081[76] << 81) +
      (src081[77] << 81) +
      (src081[78] << 81) +
      (src081[79] << 81) +
      (src081[80] << 81) +
      (src081[81] << 81) +
      (src081[82] << 81) +
      (src081[83] << 81) +
      (src081[84] << 81) +
      (src081[85] << 81) +
      (src081[86] << 81) +
      (src081[87] << 81) +
      (src081[88] << 81) +
      (src081[89] << 81) +
      (src081[90] << 81) +
      (src081[91] << 81) +
      (src081[92] << 81) +
      (src081[93] << 81) +
      (src081[94] << 81) +
      (src081[95] << 81) +
      (src081[96] << 81) +
      (src081[97] << 81) +
      (src081[98] << 81) +
      (src081[99] << 81) +
      (src081[100] << 81) +
      (src081[101] << 81) +
      (src081[102] << 81) +
      (src081[103] << 81) +
      (src081[104] << 81) +
      (src081[105] << 81) +
      (src081[106] << 81) +
      (src081[107] << 81) +
      (src081[108] << 81) +
      (src081[109] << 81) +
      (src081[110] << 81) +
      (src081[111] << 81) +
      (src081[112] << 81) +
      (src081[113] << 81) +
      (src081[114] << 81) +
      (src081[115] << 81) +
      (src081[116] << 81) +
      (src081[117] << 81) +
      (src081[118] << 81) +
      (src081[119] << 81) +
      (src081[120] << 81) +
      (src081[121] << 81) +
      (src081[122] << 81) +
      (src081[123] << 81) +
      (src081[124] << 81) +
      (src081[125] << 81) +
      (src081[126] << 81) +
      (src081[127] << 81) +
      (src082[0] << 82) +
      (src082[1] << 82) +
      (src082[2] << 82) +
      (src082[3] << 82) +
      (src082[4] << 82) +
      (src082[5] << 82) +
      (src082[6] << 82) +
      (src082[7] << 82) +
      (src082[8] << 82) +
      (src082[9] << 82) +
      (src082[10] << 82) +
      (src082[11] << 82) +
      (src082[12] << 82) +
      (src082[13] << 82) +
      (src082[14] << 82) +
      (src082[15] << 82) +
      (src082[16] << 82) +
      (src082[17] << 82) +
      (src082[18] << 82) +
      (src082[19] << 82) +
      (src082[20] << 82) +
      (src082[21] << 82) +
      (src082[22] << 82) +
      (src082[23] << 82) +
      (src082[24] << 82) +
      (src082[25] << 82) +
      (src082[26] << 82) +
      (src082[27] << 82) +
      (src082[28] << 82) +
      (src082[29] << 82) +
      (src082[30] << 82) +
      (src082[31] << 82) +
      (src082[32] << 82) +
      (src082[33] << 82) +
      (src082[34] << 82) +
      (src082[35] << 82) +
      (src082[36] << 82) +
      (src082[37] << 82) +
      (src082[38] << 82) +
      (src082[39] << 82) +
      (src082[40] << 82) +
      (src082[41] << 82) +
      (src082[42] << 82) +
      (src082[43] << 82) +
      (src082[44] << 82) +
      (src082[45] << 82) +
      (src082[46] << 82) +
      (src082[47] << 82) +
      (src082[48] << 82) +
      (src082[49] << 82) +
      (src082[50] << 82) +
      (src082[51] << 82) +
      (src082[52] << 82) +
      (src082[53] << 82) +
      (src082[54] << 82) +
      (src082[55] << 82) +
      (src082[56] << 82) +
      (src082[57] << 82) +
      (src082[58] << 82) +
      (src082[59] << 82) +
      (src082[60] << 82) +
      (src082[61] << 82) +
      (src082[62] << 82) +
      (src082[63] << 82) +
      (src082[64] << 82) +
      (src082[65] << 82) +
      (src082[66] << 82) +
      (src082[67] << 82) +
      (src082[68] << 82) +
      (src082[69] << 82) +
      (src082[70] << 82) +
      (src082[71] << 82) +
      (src082[72] << 82) +
      (src082[73] << 82) +
      (src082[74] << 82) +
      (src082[75] << 82) +
      (src082[76] << 82) +
      (src082[77] << 82) +
      (src082[78] << 82) +
      (src082[79] << 82) +
      (src082[80] << 82) +
      (src082[81] << 82) +
      (src082[82] << 82) +
      (src082[83] << 82) +
      (src082[84] << 82) +
      (src082[85] << 82) +
      (src082[86] << 82) +
      (src082[87] << 82) +
      (src082[88] << 82) +
      (src082[89] << 82) +
      (src082[90] << 82) +
      (src082[91] << 82) +
      (src082[92] << 82) +
      (src082[93] << 82) +
      (src082[94] << 82) +
      (src082[95] << 82) +
      (src082[96] << 82) +
      (src082[97] << 82) +
      (src082[98] << 82) +
      (src082[99] << 82) +
      (src082[100] << 82) +
      (src082[101] << 82) +
      (src082[102] << 82) +
      (src082[103] << 82) +
      (src082[104] << 82) +
      (src082[105] << 82) +
      (src082[106] << 82) +
      (src082[107] << 82) +
      (src082[108] << 82) +
      (src082[109] << 82) +
      (src082[110] << 82) +
      (src082[111] << 82) +
      (src082[112] << 82) +
      (src082[113] << 82) +
      (src082[114] << 82) +
      (src082[115] << 82) +
      (src082[116] << 82) +
      (src082[117] << 82) +
      (src082[118] << 82) +
      (src082[119] << 82) +
      (src082[120] << 82) +
      (src082[121] << 82) +
      (src082[122] << 82) +
      (src082[123] << 82) +
      (src082[124] << 82) +
      (src082[125] << 82) +
      (src082[126] << 82) +
      (src082[127] << 82) +
      (src083[0] << 83) +
      (src083[1] << 83) +
      (src083[2] << 83) +
      (src083[3] << 83) +
      (src083[4] << 83) +
      (src083[5] << 83) +
      (src083[6] << 83) +
      (src083[7] << 83) +
      (src083[8] << 83) +
      (src083[9] << 83) +
      (src083[10] << 83) +
      (src083[11] << 83) +
      (src083[12] << 83) +
      (src083[13] << 83) +
      (src083[14] << 83) +
      (src083[15] << 83) +
      (src083[16] << 83) +
      (src083[17] << 83) +
      (src083[18] << 83) +
      (src083[19] << 83) +
      (src083[20] << 83) +
      (src083[21] << 83) +
      (src083[22] << 83) +
      (src083[23] << 83) +
      (src083[24] << 83) +
      (src083[25] << 83) +
      (src083[26] << 83) +
      (src083[27] << 83) +
      (src083[28] << 83) +
      (src083[29] << 83) +
      (src083[30] << 83) +
      (src083[31] << 83) +
      (src083[32] << 83) +
      (src083[33] << 83) +
      (src083[34] << 83) +
      (src083[35] << 83) +
      (src083[36] << 83) +
      (src083[37] << 83) +
      (src083[38] << 83) +
      (src083[39] << 83) +
      (src083[40] << 83) +
      (src083[41] << 83) +
      (src083[42] << 83) +
      (src083[43] << 83) +
      (src083[44] << 83) +
      (src083[45] << 83) +
      (src083[46] << 83) +
      (src083[47] << 83) +
      (src083[48] << 83) +
      (src083[49] << 83) +
      (src083[50] << 83) +
      (src083[51] << 83) +
      (src083[52] << 83) +
      (src083[53] << 83) +
      (src083[54] << 83) +
      (src083[55] << 83) +
      (src083[56] << 83) +
      (src083[57] << 83) +
      (src083[58] << 83) +
      (src083[59] << 83) +
      (src083[60] << 83) +
      (src083[61] << 83) +
      (src083[62] << 83) +
      (src083[63] << 83) +
      (src083[64] << 83) +
      (src083[65] << 83) +
      (src083[66] << 83) +
      (src083[67] << 83) +
      (src083[68] << 83) +
      (src083[69] << 83) +
      (src083[70] << 83) +
      (src083[71] << 83) +
      (src083[72] << 83) +
      (src083[73] << 83) +
      (src083[74] << 83) +
      (src083[75] << 83) +
      (src083[76] << 83) +
      (src083[77] << 83) +
      (src083[78] << 83) +
      (src083[79] << 83) +
      (src083[80] << 83) +
      (src083[81] << 83) +
      (src083[82] << 83) +
      (src083[83] << 83) +
      (src083[84] << 83) +
      (src083[85] << 83) +
      (src083[86] << 83) +
      (src083[87] << 83) +
      (src083[88] << 83) +
      (src083[89] << 83) +
      (src083[90] << 83) +
      (src083[91] << 83) +
      (src083[92] << 83) +
      (src083[93] << 83) +
      (src083[94] << 83) +
      (src083[95] << 83) +
      (src083[96] << 83) +
      (src083[97] << 83) +
      (src083[98] << 83) +
      (src083[99] << 83) +
      (src083[100] << 83) +
      (src083[101] << 83) +
      (src083[102] << 83) +
      (src083[103] << 83) +
      (src083[104] << 83) +
      (src083[105] << 83) +
      (src083[106] << 83) +
      (src083[107] << 83) +
      (src083[108] << 83) +
      (src083[109] << 83) +
      (src083[110] << 83) +
      (src083[111] << 83) +
      (src083[112] << 83) +
      (src083[113] << 83) +
      (src083[114] << 83) +
      (src083[115] << 83) +
      (src083[116] << 83) +
      (src083[117] << 83) +
      (src083[118] << 83) +
      (src083[119] << 83) +
      (src083[120] << 83) +
      (src083[121] << 83) +
      (src083[122] << 83) +
      (src083[123] << 83) +
      (src083[124] << 83) +
      (src083[125] << 83) +
      (src083[126] << 83) +
      (src083[127] << 83) +
      (src084[0] << 84) +
      (src084[1] << 84) +
      (src084[2] << 84) +
      (src084[3] << 84) +
      (src084[4] << 84) +
      (src084[5] << 84) +
      (src084[6] << 84) +
      (src084[7] << 84) +
      (src084[8] << 84) +
      (src084[9] << 84) +
      (src084[10] << 84) +
      (src084[11] << 84) +
      (src084[12] << 84) +
      (src084[13] << 84) +
      (src084[14] << 84) +
      (src084[15] << 84) +
      (src084[16] << 84) +
      (src084[17] << 84) +
      (src084[18] << 84) +
      (src084[19] << 84) +
      (src084[20] << 84) +
      (src084[21] << 84) +
      (src084[22] << 84) +
      (src084[23] << 84) +
      (src084[24] << 84) +
      (src084[25] << 84) +
      (src084[26] << 84) +
      (src084[27] << 84) +
      (src084[28] << 84) +
      (src084[29] << 84) +
      (src084[30] << 84) +
      (src084[31] << 84) +
      (src084[32] << 84) +
      (src084[33] << 84) +
      (src084[34] << 84) +
      (src084[35] << 84) +
      (src084[36] << 84) +
      (src084[37] << 84) +
      (src084[38] << 84) +
      (src084[39] << 84) +
      (src084[40] << 84) +
      (src084[41] << 84) +
      (src084[42] << 84) +
      (src084[43] << 84) +
      (src084[44] << 84) +
      (src084[45] << 84) +
      (src084[46] << 84) +
      (src084[47] << 84) +
      (src084[48] << 84) +
      (src084[49] << 84) +
      (src084[50] << 84) +
      (src084[51] << 84) +
      (src084[52] << 84) +
      (src084[53] << 84) +
      (src084[54] << 84) +
      (src084[55] << 84) +
      (src084[56] << 84) +
      (src084[57] << 84) +
      (src084[58] << 84) +
      (src084[59] << 84) +
      (src084[60] << 84) +
      (src084[61] << 84) +
      (src084[62] << 84) +
      (src084[63] << 84) +
      (src084[64] << 84) +
      (src084[65] << 84) +
      (src084[66] << 84) +
      (src084[67] << 84) +
      (src084[68] << 84) +
      (src084[69] << 84) +
      (src084[70] << 84) +
      (src084[71] << 84) +
      (src084[72] << 84) +
      (src084[73] << 84) +
      (src084[74] << 84) +
      (src084[75] << 84) +
      (src084[76] << 84) +
      (src084[77] << 84) +
      (src084[78] << 84) +
      (src084[79] << 84) +
      (src084[80] << 84) +
      (src084[81] << 84) +
      (src084[82] << 84) +
      (src084[83] << 84) +
      (src084[84] << 84) +
      (src084[85] << 84) +
      (src084[86] << 84) +
      (src084[87] << 84) +
      (src084[88] << 84) +
      (src084[89] << 84) +
      (src084[90] << 84) +
      (src084[91] << 84) +
      (src084[92] << 84) +
      (src084[93] << 84) +
      (src084[94] << 84) +
      (src084[95] << 84) +
      (src084[96] << 84) +
      (src084[97] << 84) +
      (src084[98] << 84) +
      (src084[99] << 84) +
      (src084[100] << 84) +
      (src084[101] << 84) +
      (src084[102] << 84) +
      (src084[103] << 84) +
      (src084[104] << 84) +
      (src084[105] << 84) +
      (src084[106] << 84) +
      (src084[107] << 84) +
      (src084[108] << 84) +
      (src084[109] << 84) +
      (src084[110] << 84) +
      (src084[111] << 84) +
      (src084[112] << 84) +
      (src084[113] << 84) +
      (src084[114] << 84) +
      (src084[115] << 84) +
      (src084[116] << 84) +
      (src084[117] << 84) +
      (src084[118] << 84) +
      (src084[119] << 84) +
      (src084[120] << 84) +
      (src084[121] << 84) +
      (src084[122] << 84) +
      (src084[123] << 84) +
      (src084[124] << 84) +
      (src084[125] << 84) +
      (src084[126] << 84) +
      (src084[127] << 84) +
      (src085[0] << 85) +
      (src085[1] << 85) +
      (src085[2] << 85) +
      (src085[3] << 85) +
      (src085[4] << 85) +
      (src085[5] << 85) +
      (src085[6] << 85) +
      (src085[7] << 85) +
      (src085[8] << 85) +
      (src085[9] << 85) +
      (src085[10] << 85) +
      (src085[11] << 85) +
      (src085[12] << 85) +
      (src085[13] << 85) +
      (src085[14] << 85) +
      (src085[15] << 85) +
      (src085[16] << 85) +
      (src085[17] << 85) +
      (src085[18] << 85) +
      (src085[19] << 85) +
      (src085[20] << 85) +
      (src085[21] << 85) +
      (src085[22] << 85) +
      (src085[23] << 85) +
      (src085[24] << 85) +
      (src085[25] << 85) +
      (src085[26] << 85) +
      (src085[27] << 85) +
      (src085[28] << 85) +
      (src085[29] << 85) +
      (src085[30] << 85) +
      (src085[31] << 85) +
      (src085[32] << 85) +
      (src085[33] << 85) +
      (src085[34] << 85) +
      (src085[35] << 85) +
      (src085[36] << 85) +
      (src085[37] << 85) +
      (src085[38] << 85) +
      (src085[39] << 85) +
      (src085[40] << 85) +
      (src085[41] << 85) +
      (src085[42] << 85) +
      (src085[43] << 85) +
      (src085[44] << 85) +
      (src085[45] << 85) +
      (src085[46] << 85) +
      (src085[47] << 85) +
      (src085[48] << 85) +
      (src085[49] << 85) +
      (src085[50] << 85) +
      (src085[51] << 85) +
      (src085[52] << 85) +
      (src085[53] << 85) +
      (src085[54] << 85) +
      (src085[55] << 85) +
      (src085[56] << 85) +
      (src085[57] << 85) +
      (src085[58] << 85) +
      (src085[59] << 85) +
      (src085[60] << 85) +
      (src085[61] << 85) +
      (src085[62] << 85) +
      (src085[63] << 85) +
      (src085[64] << 85) +
      (src085[65] << 85) +
      (src085[66] << 85) +
      (src085[67] << 85) +
      (src085[68] << 85) +
      (src085[69] << 85) +
      (src085[70] << 85) +
      (src085[71] << 85) +
      (src085[72] << 85) +
      (src085[73] << 85) +
      (src085[74] << 85) +
      (src085[75] << 85) +
      (src085[76] << 85) +
      (src085[77] << 85) +
      (src085[78] << 85) +
      (src085[79] << 85) +
      (src085[80] << 85) +
      (src085[81] << 85) +
      (src085[82] << 85) +
      (src085[83] << 85) +
      (src085[84] << 85) +
      (src085[85] << 85) +
      (src085[86] << 85) +
      (src085[87] << 85) +
      (src085[88] << 85) +
      (src085[89] << 85) +
      (src085[90] << 85) +
      (src085[91] << 85) +
      (src085[92] << 85) +
      (src085[93] << 85) +
      (src085[94] << 85) +
      (src085[95] << 85) +
      (src085[96] << 85) +
      (src085[97] << 85) +
      (src085[98] << 85) +
      (src085[99] << 85) +
      (src085[100] << 85) +
      (src085[101] << 85) +
      (src085[102] << 85) +
      (src085[103] << 85) +
      (src085[104] << 85) +
      (src085[105] << 85) +
      (src085[106] << 85) +
      (src085[107] << 85) +
      (src085[108] << 85) +
      (src085[109] << 85) +
      (src085[110] << 85) +
      (src085[111] << 85) +
      (src085[112] << 85) +
      (src085[113] << 85) +
      (src085[114] << 85) +
      (src085[115] << 85) +
      (src085[116] << 85) +
      (src085[117] << 85) +
      (src085[118] << 85) +
      (src085[119] << 85) +
      (src085[120] << 85) +
      (src085[121] << 85) +
      (src085[122] << 85) +
      (src085[123] << 85) +
      (src085[124] << 85) +
      (src085[125] << 85) +
      (src085[126] << 85) +
      (src085[127] << 85) +
      (src086[0] << 86) +
      (src086[1] << 86) +
      (src086[2] << 86) +
      (src086[3] << 86) +
      (src086[4] << 86) +
      (src086[5] << 86) +
      (src086[6] << 86) +
      (src086[7] << 86) +
      (src086[8] << 86) +
      (src086[9] << 86) +
      (src086[10] << 86) +
      (src086[11] << 86) +
      (src086[12] << 86) +
      (src086[13] << 86) +
      (src086[14] << 86) +
      (src086[15] << 86) +
      (src086[16] << 86) +
      (src086[17] << 86) +
      (src086[18] << 86) +
      (src086[19] << 86) +
      (src086[20] << 86) +
      (src086[21] << 86) +
      (src086[22] << 86) +
      (src086[23] << 86) +
      (src086[24] << 86) +
      (src086[25] << 86) +
      (src086[26] << 86) +
      (src086[27] << 86) +
      (src086[28] << 86) +
      (src086[29] << 86) +
      (src086[30] << 86) +
      (src086[31] << 86) +
      (src086[32] << 86) +
      (src086[33] << 86) +
      (src086[34] << 86) +
      (src086[35] << 86) +
      (src086[36] << 86) +
      (src086[37] << 86) +
      (src086[38] << 86) +
      (src086[39] << 86) +
      (src086[40] << 86) +
      (src086[41] << 86) +
      (src086[42] << 86) +
      (src086[43] << 86) +
      (src086[44] << 86) +
      (src086[45] << 86) +
      (src086[46] << 86) +
      (src086[47] << 86) +
      (src086[48] << 86) +
      (src086[49] << 86) +
      (src086[50] << 86) +
      (src086[51] << 86) +
      (src086[52] << 86) +
      (src086[53] << 86) +
      (src086[54] << 86) +
      (src086[55] << 86) +
      (src086[56] << 86) +
      (src086[57] << 86) +
      (src086[58] << 86) +
      (src086[59] << 86) +
      (src086[60] << 86) +
      (src086[61] << 86) +
      (src086[62] << 86) +
      (src086[63] << 86) +
      (src086[64] << 86) +
      (src086[65] << 86) +
      (src086[66] << 86) +
      (src086[67] << 86) +
      (src086[68] << 86) +
      (src086[69] << 86) +
      (src086[70] << 86) +
      (src086[71] << 86) +
      (src086[72] << 86) +
      (src086[73] << 86) +
      (src086[74] << 86) +
      (src086[75] << 86) +
      (src086[76] << 86) +
      (src086[77] << 86) +
      (src086[78] << 86) +
      (src086[79] << 86) +
      (src086[80] << 86) +
      (src086[81] << 86) +
      (src086[82] << 86) +
      (src086[83] << 86) +
      (src086[84] << 86) +
      (src086[85] << 86) +
      (src086[86] << 86) +
      (src086[87] << 86) +
      (src086[88] << 86) +
      (src086[89] << 86) +
      (src086[90] << 86) +
      (src086[91] << 86) +
      (src086[92] << 86) +
      (src086[93] << 86) +
      (src086[94] << 86) +
      (src086[95] << 86) +
      (src086[96] << 86) +
      (src086[97] << 86) +
      (src086[98] << 86) +
      (src086[99] << 86) +
      (src086[100] << 86) +
      (src086[101] << 86) +
      (src086[102] << 86) +
      (src086[103] << 86) +
      (src086[104] << 86) +
      (src086[105] << 86) +
      (src086[106] << 86) +
      (src086[107] << 86) +
      (src086[108] << 86) +
      (src086[109] << 86) +
      (src086[110] << 86) +
      (src086[111] << 86) +
      (src086[112] << 86) +
      (src086[113] << 86) +
      (src086[114] << 86) +
      (src086[115] << 86) +
      (src086[116] << 86) +
      (src086[117] << 86) +
      (src086[118] << 86) +
      (src086[119] << 86) +
      (src086[120] << 86) +
      (src086[121] << 86) +
      (src086[122] << 86) +
      (src086[123] << 86) +
      (src086[124] << 86) +
      (src086[125] << 86) +
      (src086[126] << 86) +
      (src086[127] << 86) +
      (src087[0] << 87) +
      (src087[1] << 87) +
      (src087[2] << 87) +
      (src087[3] << 87) +
      (src087[4] << 87) +
      (src087[5] << 87) +
      (src087[6] << 87) +
      (src087[7] << 87) +
      (src087[8] << 87) +
      (src087[9] << 87) +
      (src087[10] << 87) +
      (src087[11] << 87) +
      (src087[12] << 87) +
      (src087[13] << 87) +
      (src087[14] << 87) +
      (src087[15] << 87) +
      (src087[16] << 87) +
      (src087[17] << 87) +
      (src087[18] << 87) +
      (src087[19] << 87) +
      (src087[20] << 87) +
      (src087[21] << 87) +
      (src087[22] << 87) +
      (src087[23] << 87) +
      (src087[24] << 87) +
      (src087[25] << 87) +
      (src087[26] << 87) +
      (src087[27] << 87) +
      (src087[28] << 87) +
      (src087[29] << 87) +
      (src087[30] << 87) +
      (src087[31] << 87) +
      (src087[32] << 87) +
      (src087[33] << 87) +
      (src087[34] << 87) +
      (src087[35] << 87) +
      (src087[36] << 87) +
      (src087[37] << 87) +
      (src087[38] << 87) +
      (src087[39] << 87) +
      (src087[40] << 87) +
      (src087[41] << 87) +
      (src087[42] << 87) +
      (src087[43] << 87) +
      (src087[44] << 87) +
      (src087[45] << 87) +
      (src087[46] << 87) +
      (src087[47] << 87) +
      (src087[48] << 87) +
      (src087[49] << 87) +
      (src087[50] << 87) +
      (src087[51] << 87) +
      (src087[52] << 87) +
      (src087[53] << 87) +
      (src087[54] << 87) +
      (src087[55] << 87) +
      (src087[56] << 87) +
      (src087[57] << 87) +
      (src087[58] << 87) +
      (src087[59] << 87) +
      (src087[60] << 87) +
      (src087[61] << 87) +
      (src087[62] << 87) +
      (src087[63] << 87) +
      (src087[64] << 87) +
      (src087[65] << 87) +
      (src087[66] << 87) +
      (src087[67] << 87) +
      (src087[68] << 87) +
      (src087[69] << 87) +
      (src087[70] << 87) +
      (src087[71] << 87) +
      (src087[72] << 87) +
      (src087[73] << 87) +
      (src087[74] << 87) +
      (src087[75] << 87) +
      (src087[76] << 87) +
      (src087[77] << 87) +
      (src087[78] << 87) +
      (src087[79] << 87) +
      (src087[80] << 87) +
      (src087[81] << 87) +
      (src087[82] << 87) +
      (src087[83] << 87) +
      (src087[84] << 87) +
      (src087[85] << 87) +
      (src087[86] << 87) +
      (src087[87] << 87) +
      (src087[88] << 87) +
      (src087[89] << 87) +
      (src087[90] << 87) +
      (src087[91] << 87) +
      (src087[92] << 87) +
      (src087[93] << 87) +
      (src087[94] << 87) +
      (src087[95] << 87) +
      (src087[96] << 87) +
      (src087[97] << 87) +
      (src087[98] << 87) +
      (src087[99] << 87) +
      (src087[100] << 87) +
      (src087[101] << 87) +
      (src087[102] << 87) +
      (src087[103] << 87) +
      (src087[104] << 87) +
      (src087[105] << 87) +
      (src087[106] << 87) +
      (src087[107] << 87) +
      (src087[108] << 87) +
      (src087[109] << 87) +
      (src087[110] << 87) +
      (src087[111] << 87) +
      (src087[112] << 87) +
      (src087[113] << 87) +
      (src087[114] << 87) +
      (src087[115] << 87) +
      (src087[116] << 87) +
      (src087[117] << 87) +
      (src087[118] << 87) +
      (src087[119] << 87) +
      (src087[120] << 87) +
      (src087[121] << 87) +
      (src087[122] << 87) +
      (src087[123] << 87) +
      (src087[124] << 87) +
      (src087[125] << 87) +
      (src087[126] << 87) +
      (src087[127] << 87) +
      (src088[0] << 88) +
      (src088[1] << 88) +
      (src088[2] << 88) +
      (src088[3] << 88) +
      (src088[4] << 88) +
      (src088[5] << 88) +
      (src088[6] << 88) +
      (src088[7] << 88) +
      (src088[8] << 88) +
      (src088[9] << 88) +
      (src088[10] << 88) +
      (src088[11] << 88) +
      (src088[12] << 88) +
      (src088[13] << 88) +
      (src088[14] << 88) +
      (src088[15] << 88) +
      (src088[16] << 88) +
      (src088[17] << 88) +
      (src088[18] << 88) +
      (src088[19] << 88) +
      (src088[20] << 88) +
      (src088[21] << 88) +
      (src088[22] << 88) +
      (src088[23] << 88) +
      (src088[24] << 88) +
      (src088[25] << 88) +
      (src088[26] << 88) +
      (src088[27] << 88) +
      (src088[28] << 88) +
      (src088[29] << 88) +
      (src088[30] << 88) +
      (src088[31] << 88) +
      (src088[32] << 88) +
      (src088[33] << 88) +
      (src088[34] << 88) +
      (src088[35] << 88) +
      (src088[36] << 88) +
      (src088[37] << 88) +
      (src088[38] << 88) +
      (src088[39] << 88) +
      (src088[40] << 88) +
      (src088[41] << 88) +
      (src088[42] << 88) +
      (src088[43] << 88) +
      (src088[44] << 88) +
      (src088[45] << 88) +
      (src088[46] << 88) +
      (src088[47] << 88) +
      (src088[48] << 88) +
      (src088[49] << 88) +
      (src088[50] << 88) +
      (src088[51] << 88) +
      (src088[52] << 88) +
      (src088[53] << 88) +
      (src088[54] << 88) +
      (src088[55] << 88) +
      (src088[56] << 88) +
      (src088[57] << 88) +
      (src088[58] << 88) +
      (src088[59] << 88) +
      (src088[60] << 88) +
      (src088[61] << 88) +
      (src088[62] << 88) +
      (src088[63] << 88) +
      (src088[64] << 88) +
      (src088[65] << 88) +
      (src088[66] << 88) +
      (src088[67] << 88) +
      (src088[68] << 88) +
      (src088[69] << 88) +
      (src088[70] << 88) +
      (src088[71] << 88) +
      (src088[72] << 88) +
      (src088[73] << 88) +
      (src088[74] << 88) +
      (src088[75] << 88) +
      (src088[76] << 88) +
      (src088[77] << 88) +
      (src088[78] << 88) +
      (src088[79] << 88) +
      (src088[80] << 88) +
      (src088[81] << 88) +
      (src088[82] << 88) +
      (src088[83] << 88) +
      (src088[84] << 88) +
      (src088[85] << 88) +
      (src088[86] << 88) +
      (src088[87] << 88) +
      (src088[88] << 88) +
      (src088[89] << 88) +
      (src088[90] << 88) +
      (src088[91] << 88) +
      (src088[92] << 88) +
      (src088[93] << 88) +
      (src088[94] << 88) +
      (src088[95] << 88) +
      (src088[96] << 88) +
      (src088[97] << 88) +
      (src088[98] << 88) +
      (src088[99] << 88) +
      (src088[100] << 88) +
      (src088[101] << 88) +
      (src088[102] << 88) +
      (src088[103] << 88) +
      (src088[104] << 88) +
      (src088[105] << 88) +
      (src088[106] << 88) +
      (src088[107] << 88) +
      (src088[108] << 88) +
      (src088[109] << 88) +
      (src088[110] << 88) +
      (src088[111] << 88) +
      (src088[112] << 88) +
      (src088[113] << 88) +
      (src088[114] << 88) +
      (src088[115] << 88) +
      (src088[116] << 88) +
      (src088[117] << 88) +
      (src088[118] << 88) +
      (src088[119] << 88) +
      (src088[120] << 88) +
      (src088[121] << 88) +
      (src088[122] << 88) +
      (src088[123] << 88) +
      (src088[124] << 88) +
      (src088[125] << 88) +
      (src088[126] << 88) +
      (src088[127] << 88) +
      (src089[0] << 89) +
      (src089[1] << 89) +
      (src089[2] << 89) +
      (src089[3] << 89) +
      (src089[4] << 89) +
      (src089[5] << 89) +
      (src089[6] << 89) +
      (src089[7] << 89) +
      (src089[8] << 89) +
      (src089[9] << 89) +
      (src089[10] << 89) +
      (src089[11] << 89) +
      (src089[12] << 89) +
      (src089[13] << 89) +
      (src089[14] << 89) +
      (src089[15] << 89) +
      (src089[16] << 89) +
      (src089[17] << 89) +
      (src089[18] << 89) +
      (src089[19] << 89) +
      (src089[20] << 89) +
      (src089[21] << 89) +
      (src089[22] << 89) +
      (src089[23] << 89) +
      (src089[24] << 89) +
      (src089[25] << 89) +
      (src089[26] << 89) +
      (src089[27] << 89) +
      (src089[28] << 89) +
      (src089[29] << 89) +
      (src089[30] << 89) +
      (src089[31] << 89) +
      (src089[32] << 89) +
      (src089[33] << 89) +
      (src089[34] << 89) +
      (src089[35] << 89) +
      (src089[36] << 89) +
      (src089[37] << 89) +
      (src089[38] << 89) +
      (src089[39] << 89) +
      (src089[40] << 89) +
      (src089[41] << 89) +
      (src089[42] << 89) +
      (src089[43] << 89) +
      (src089[44] << 89) +
      (src089[45] << 89) +
      (src089[46] << 89) +
      (src089[47] << 89) +
      (src089[48] << 89) +
      (src089[49] << 89) +
      (src089[50] << 89) +
      (src089[51] << 89) +
      (src089[52] << 89) +
      (src089[53] << 89) +
      (src089[54] << 89) +
      (src089[55] << 89) +
      (src089[56] << 89) +
      (src089[57] << 89) +
      (src089[58] << 89) +
      (src089[59] << 89) +
      (src089[60] << 89) +
      (src089[61] << 89) +
      (src089[62] << 89) +
      (src089[63] << 89) +
      (src089[64] << 89) +
      (src089[65] << 89) +
      (src089[66] << 89) +
      (src089[67] << 89) +
      (src089[68] << 89) +
      (src089[69] << 89) +
      (src089[70] << 89) +
      (src089[71] << 89) +
      (src089[72] << 89) +
      (src089[73] << 89) +
      (src089[74] << 89) +
      (src089[75] << 89) +
      (src089[76] << 89) +
      (src089[77] << 89) +
      (src089[78] << 89) +
      (src089[79] << 89) +
      (src089[80] << 89) +
      (src089[81] << 89) +
      (src089[82] << 89) +
      (src089[83] << 89) +
      (src089[84] << 89) +
      (src089[85] << 89) +
      (src089[86] << 89) +
      (src089[87] << 89) +
      (src089[88] << 89) +
      (src089[89] << 89) +
      (src089[90] << 89) +
      (src089[91] << 89) +
      (src089[92] << 89) +
      (src089[93] << 89) +
      (src089[94] << 89) +
      (src089[95] << 89) +
      (src089[96] << 89) +
      (src089[97] << 89) +
      (src089[98] << 89) +
      (src089[99] << 89) +
      (src089[100] << 89) +
      (src089[101] << 89) +
      (src089[102] << 89) +
      (src089[103] << 89) +
      (src089[104] << 89) +
      (src089[105] << 89) +
      (src089[106] << 89) +
      (src089[107] << 89) +
      (src089[108] << 89) +
      (src089[109] << 89) +
      (src089[110] << 89) +
      (src089[111] << 89) +
      (src089[112] << 89) +
      (src089[113] << 89) +
      (src089[114] << 89) +
      (src089[115] << 89) +
      (src089[116] << 89) +
      (src089[117] << 89) +
      (src089[118] << 89) +
      (src089[119] << 89) +
      (src089[120] << 89) +
      (src089[121] << 89) +
      (src089[122] << 89) +
      (src089[123] << 89) +
      (src089[124] << 89) +
      (src089[125] << 89) +
      (src089[126] << 89) +
      (src089[127] << 89) +
      (src090[0] << 90) +
      (src090[1] << 90) +
      (src090[2] << 90) +
      (src090[3] << 90) +
      (src090[4] << 90) +
      (src090[5] << 90) +
      (src090[6] << 90) +
      (src090[7] << 90) +
      (src090[8] << 90) +
      (src090[9] << 90) +
      (src090[10] << 90) +
      (src090[11] << 90) +
      (src090[12] << 90) +
      (src090[13] << 90) +
      (src090[14] << 90) +
      (src090[15] << 90) +
      (src090[16] << 90) +
      (src090[17] << 90) +
      (src090[18] << 90) +
      (src090[19] << 90) +
      (src090[20] << 90) +
      (src090[21] << 90) +
      (src090[22] << 90) +
      (src090[23] << 90) +
      (src090[24] << 90) +
      (src090[25] << 90) +
      (src090[26] << 90) +
      (src090[27] << 90) +
      (src090[28] << 90) +
      (src090[29] << 90) +
      (src090[30] << 90) +
      (src090[31] << 90) +
      (src090[32] << 90) +
      (src090[33] << 90) +
      (src090[34] << 90) +
      (src090[35] << 90) +
      (src090[36] << 90) +
      (src090[37] << 90) +
      (src090[38] << 90) +
      (src090[39] << 90) +
      (src090[40] << 90) +
      (src090[41] << 90) +
      (src090[42] << 90) +
      (src090[43] << 90) +
      (src090[44] << 90) +
      (src090[45] << 90) +
      (src090[46] << 90) +
      (src090[47] << 90) +
      (src090[48] << 90) +
      (src090[49] << 90) +
      (src090[50] << 90) +
      (src090[51] << 90) +
      (src090[52] << 90) +
      (src090[53] << 90) +
      (src090[54] << 90) +
      (src090[55] << 90) +
      (src090[56] << 90) +
      (src090[57] << 90) +
      (src090[58] << 90) +
      (src090[59] << 90) +
      (src090[60] << 90) +
      (src090[61] << 90) +
      (src090[62] << 90) +
      (src090[63] << 90) +
      (src090[64] << 90) +
      (src090[65] << 90) +
      (src090[66] << 90) +
      (src090[67] << 90) +
      (src090[68] << 90) +
      (src090[69] << 90) +
      (src090[70] << 90) +
      (src090[71] << 90) +
      (src090[72] << 90) +
      (src090[73] << 90) +
      (src090[74] << 90) +
      (src090[75] << 90) +
      (src090[76] << 90) +
      (src090[77] << 90) +
      (src090[78] << 90) +
      (src090[79] << 90) +
      (src090[80] << 90) +
      (src090[81] << 90) +
      (src090[82] << 90) +
      (src090[83] << 90) +
      (src090[84] << 90) +
      (src090[85] << 90) +
      (src090[86] << 90) +
      (src090[87] << 90) +
      (src090[88] << 90) +
      (src090[89] << 90) +
      (src090[90] << 90) +
      (src090[91] << 90) +
      (src090[92] << 90) +
      (src090[93] << 90) +
      (src090[94] << 90) +
      (src090[95] << 90) +
      (src090[96] << 90) +
      (src090[97] << 90) +
      (src090[98] << 90) +
      (src090[99] << 90) +
      (src090[100] << 90) +
      (src090[101] << 90) +
      (src090[102] << 90) +
      (src090[103] << 90) +
      (src090[104] << 90) +
      (src090[105] << 90) +
      (src090[106] << 90) +
      (src090[107] << 90) +
      (src090[108] << 90) +
      (src090[109] << 90) +
      (src090[110] << 90) +
      (src090[111] << 90) +
      (src090[112] << 90) +
      (src090[113] << 90) +
      (src090[114] << 90) +
      (src090[115] << 90) +
      (src090[116] << 90) +
      (src090[117] << 90) +
      (src090[118] << 90) +
      (src090[119] << 90) +
      (src090[120] << 90) +
      (src090[121] << 90) +
      (src090[122] << 90) +
      (src090[123] << 90) +
      (src090[124] << 90) +
      (src090[125] << 90) +
      (src090[126] << 90) +
      (src090[127] << 90) +
      (src091[0] << 91) +
      (src091[1] << 91) +
      (src091[2] << 91) +
      (src091[3] << 91) +
      (src091[4] << 91) +
      (src091[5] << 91) +
      (src091[6] << 91) +
      (src091[7] << 91) +
      (src091[8] << 91) +
      (src091[9] << 91) +
      (src091[10] << 91) +
      (src091[11] << 91) +
      (src091[12] << 91) +
      (src091[13] << 91) +
      (src091[14] << 91) +
      (src091[15] << 91) +
      (src091[16] << 91) +
      (src091[17] << 91) +
      (src091[18] << 91) +
      (src091[19] << 91) +
      (src091[20] << 91) +
      (src091[21] << 91) +
      (src091[22] << 91) +
      (src091[23] << 91) +
      (src091[24] << 91) +
      (src091[25] << 91) +
      (src091[26] << 91) +
      (src091[27] << 91) +
      (src091[28] << 91) +
      (src091[29] << 91) +
      (src091[30] << 91) +
      (src091[31] << 91) +
      (src091[32] << 91) +
      (src091[33] << 91) +
      (src091[34] << 91) +
      (src091[35] << 91) +
      (src091[36] << 91) +
      (src091[37] << 91) +
      (src091[38] << 91) +
      (src091[39] << 91) +
      (src091[40] << 91) +
      (src091[41] << 91) +
      (src091[42] << 91) +
      (src091[43] << 91) +
      (src091[44] << 91) +
      (src091[45] << 91) +
      (src091[46] << 91) +
      (src091[47] << 91) +
      (src091[48] << 91) +
      (src091[49] << 91) +
      (src091[50] << 91) +
      (src091[51] << 91) +
      (src091[52] << 91) +
      (src091[53] << 91) +
      (src091[54] << 91) +
      (src091[55] << 91) +
      (src091[56] << 91) +
      (src091[57] << 91) +
      (src091[58] << 91) +
      (src091[59] << 91) +
      (src091[60] << 91) +
      (src091[61] << 91) +
      (src091[62] << 91) +
      (src091[63] << 91) +
      (src091[64] << 91) +
      (src091[65] << 91) +
      (src091[66] << 91) +
      (src091[67] << 91) +
      (src091[68] << 91) +
      (src091[69] << 91) +
      (src091[70] << 91) +
      (src091[71] << 91) +
      (src091[72] << 91) +
      (src091[73] << 91) +
      (src091[74] << 91) +
      (src091[75] << 91) +
      (src091[76] << 91) +
      (src091[77] << 91) +
      (src091[78] << 91) +
      (src091[79] << 91) +
      (src091[80] << 91) +
      (src091[81] << 91) +
      (src091[82] << 91) +
      (src091[83] << 91) +
      (src091[84] << 91) +
      (src091[85] << 91) +
      (src091[86] << 91) +
      (src091[87] << 91) +
      (src091[88] << 91) +
      (src091[89] << 91) +
      (src091[90] << 91) +
      (src091[91] << 91) +
      (src091[92] << 91) +
      (src091[93] << 91) +
      (src091[94] << 91) +
      (src091[95] << 91) +
      (src091[96] << 91) +
      (src091[97] << 91) +
      (src091[98] << 91) +
      (src091[99] << 91) +
      (src091[100] << 91) +
      (src091[101] << 91) +
      (src091[102] << 91) +
      (src091[103] << 91) +
      (src091[104] << 91) +
      (src091[105] << 91) +
      (src091[106] << 91) +
      (src091[107] << 91) +
      (src091[108] << 91) +
      (src091[109] << 91) +
      (src091[110] << 91) +
      (src091[111] << 91) +
      (src091[112] << 91) +
      (src091[113] << 91) +
      (src091[114] << 91) +
      (src091[115] << 91) +
      (src091[116] << 91) +
      (src091[117] << 91) +
      (src091[118] << 91) +
      (src091[119] << 91) +
      (src091[120] << 91) +
      (src091[121] << 91) +
      (src091[122] << 91) +
      (src091[123] << 91) +
      (src091[124] << 91) +
      (src091[125] << 91) +
      (src091[126] << 91) +
      (src091[127] << 91) +
      (src092[0] << 92) +
      (src092[1] << 92) +
      (src092[2] << 92) +
      (src092[3] << 92) +
      (src092[4] << 92) +
      (src092[5] << 92) +
      (src092[6] << 92) +
      (src092[7] << 92) +
      (src092[8] << 92) +
      (src092[9] << 92) +
      (src092[10] << 92) +
      (src092[11] << 92) +
      (src092[12] << 92) +
      (src092[13] << 92) +
      (src092[14] << 92) +
      (src092[15] << 92) +
      (src092[16] << 92) +
      (src092[17] << 92) +
      (src092[18] << 92) +
      (src092[19] << 92) +
      (src092[20] << 92) +
      (src092[21] << 92) +
      (src092[22] << 92) +
      (src092[23] << 92) +
      (src092[24] << 92) +
      (src092[25] << 92) +
      (src092[26] << 92) +
      (src092[27] << 92) +
      (src092[28] << 92) +
      (src092[29] << 92) +
      (src092[30] << 92) +
      (src092[31] << 92) +
      (src092[32] << 92) +
      (src092[33] << 92) +
      (src092[34] << 92) +
      (src092[35] << 92) +
      (src092[36] << 92) +
      (src092[37] << 92) +
      (src092[38] << 92) +
      (src092[39] << 92) +
      (src092[40] << 92) +
      (src092[41] << 92) +
      (src092[42] << 92) +
      (src092[43] << 92) +
      (src092[44] << 92) +
      (src092[45] << 92) +
      (src092[46] << 92) +
      (src092[47] << 92) +
      (src092[48] << 92) +
      (src092[49] << 92) +
      (src092[50] << 92) +
      (src092[51] << 92) +
      (src092[52] << 92) +
      (src092[53] << 92) +
      (src092[54] << 92) +
      (src092[55] << 92) +
      (src092[56] << 92) +
      (src092[57] << 92) +
      (src092[58] << 92) +
      (src092[59] << 92) +
      (src092[60] << 92) +
      (src092[61] << 92) +
      (src092[62] << 92) +
      (src092[63] << 92) +
      (src092[64] << 92) +
      (src092[65] << 92) +
      (src092[66] << 92) +
      (src092[67] << 92) +
      (src092[68] << 92) +
      (src092[69] << 92) +
      (src092[70] << 92) +
      (src092[71] << 92) +
      (src092[72] << 92) +
      (src092[73] << 92) +
      (src092[74] << 92) +
      (src092[75] << 92) +
      (src092[76] << 92) +
      (src092[77] << 92) +
      (src092[78] << 92) +
      (src092[79] << 92) +
      (src092[80] << 92) +
      (src092[81] << 92) +
      (src092[82] << 92) +
      (src092[83] << 92) +
      (src092[84] << 92) +
      (src092[85] << 92) +
      (src092[86] << 92) +
      (src092[87] << 92) +
      (src092[88] << 92) +
      (src092[89] << 92) +
      (src092[90] << 92) +
      (src092[91] << 92) +
      (src092[92] << 92) +
      (src092[93] << 92) +
      (src092[94] << 92) +
      (src092[95] << 92) +
      (src092[96] << 92) +
      (src092[97] << 92) +
      (src092[98] << 92) +
      (src092[99] << 92) +
      (src092[100] << 92) +
      (src092[101] << 92) +
      (src092[102] << 92) +
      (src092[103] << 92) +
      (src092[104] << 92) +
      (src092[105] << 92) +
      (src092[106] << 92) +
      (src092[107] << 92) +
      (src092[108] << 92) +
      (src092[109] << 92) +
      (src092[110] << 92) +
      (src092[111] << 92) +
      (src092[112] << 92) +
      (src092[113] << 92) +
      (src092[114] << 92) +
      (src092[115] << 92) +
      (src092[116] << 92) +
      (src092[117] << 92) +
      (src092[118] << 92) +
      (src092[119] << 92) +
      (src092[120] << 92) +
      (src092[121] << 92) +
      (src092[122] << 92) +
      (src092[123] << 92) +
      (src092[124] << 92) +
      (src092[125] << 92) +
      (src092[126] << 92) +
      (src092[127] << 92) +
      (src093[0] << 93) +
      (src093[1] << 93) +
      (src093[2] << 93) +
      (src093[3] << 93) +
      (src093[4] << 93) +
      (src093[5] << 93) +
      (src093[6] << 93) +
      (src093[7] << 93) +
      (src093[8] << 93) +
      (src093[9] << 93) +
      (src093[10] << 93) +
      (src093[11] << 93) +
      (src093[12] << 93) +
      (src093[13] << 93) +
      (src093[14] << 93) +
      (src093[15] << 93) +
      (src093[16] << 93) +
      (src093[17] << 93) +
      (src093[18] << 93) +
      (src093[19] << 93) +
      (src093[20] << 93) +
      (src093[21] << 93) +
      (src093[22] << 93) +
      (src093[23] << 93) +
      (src093[24] << 93) +
      (src093[25] << 93) +
      (src093[26] << 93) +
      (src093[27] << 93) +
      (src093[28] << 93) +
      (src093[29] << 93) +
      (src093[30] << 93) +
      (src093[31] << 93) +
      (src093[32] << 93) +
      (src093[33] << 93) +
      (src093[34] << 93) +
      (src093[35] << 93) +
      (src093[36] << 93) +
      (src093[37] << 93) +
      (src093[38] << 93) +
      (src093[39] << 93) +
      (src093[40] << 93) +
      (src093[41] << 93) +
      (src093[42] << 93) +
      (src093[43] << 93) +
      (src093[44] << 93) +
      (src093[45] << 93) +
      (src093[46] << 93) +
      (src093[47] << 93) +
      (src093[48] << 93) +
      (src093[49] << 93) +
      (src093[50] << 93) +
      (src093[51] << 93) +
      (src093[52] << 93) +
      (src093[53] << 93) +
      (src093[54] << 93) +
      (src093[55] << 93) +
      (src093[56] << 93) +
      (src093[57] << 93) +
      (src093[58] << 93) +
      (src093[59] << 93) +
      (src093[60] << 93) +
      (src093[61] << 93) +
      (src093[62] << 93) +
      (src093[63] << 93) +
      (src093[64] << 93) +
      (src093[65] << 93) +
      (src093[66] << 93) +
      (src093[67] << 93) +
      (src093[68] << 93) +
      (src093[69] << 93) +
      (src093[70] << 93) +
      (src093[71] << 93) +
      (src093[72] << 93) +
      (src093[73] << 93) +
      (src093[74] << 93) +
      (src093[75] << 93) +
      (src093[76] << 93) +
      (src093[77] << 93) +
      (src093[78] << 93) +
      (src093[79] << 93) +
      (src093[80] << 93) +
      (src093[81] << 93) +
      (src093[82] << 93) +
      (src093[83] << 93) +
      (src093[84] << 93) +
      (src093[85] << 93) +
      (src093[86] << 93) +
      (src093[87] << 93) +
      (src093[88] << 93) +
      (src093[89] << 93) +
      (src093[90] << 93) +
      (src093[91] << 93) +
      (src093[92] << 93) +
      (src093[93] << 93) +
      (src093[94] << 93) +
      (src093[95] << 93) +
      (src093[96] << 93) +
      (src093[97] << 93) +
      (src093[98] << 93) +
      (src093[99] << 93) +
      (src093[100] << 93) +
      (src093[101] << 93) +
      (src093[102] << 93) +
      (src093[103] << 93) +
      (src093[104] << 93) +
      (src093[105] << 93) +
      (src093[106] << 93) +
      (src093[107] << 93) +
      (src093[108] << 93) +
      (src093[109] << 93) +
      (src093[110] << 93) +
      (src093[111] << 93) +
      (src093[112] << 93) +
      (src093[113] << 93) +
      (src093[114] << 93) +
      (src093[115] << 93) +
      (src093[116] << 93) +
      (src093[117] << 93) +
      (src093[118] << 93) +
      (src093[119] << 93) +
      (src093[120] << 93) +
      (src093[121] << 93) +
      (src093[122] << 93) +
      (src093[123] << 93) +
      (src093[124] << 93) +
      (src093[125] << 93) +
      (src093[126] << 93) +
      (src093[127] << 93) +
      (src094[0] << 94) +
      (src094[1] << 94) +
      (src094[2] << 94) +
      (src094[3] << 94) +
      (src094[4] << 94) +
      (src094[5] << 94) +
      (src094[6] << 94) +
      (src094[7] << 94) +
      (src094[8] << 94) +
      (src094[9] << 94) +
      (src094[10] << 94) +
      (src094[11] << 94) +
      (src094[12] << 94) +
      (src094[13] << 94) +
      (src094[14] << 94) +
      (src094[15] << 94) +
      (src094[16] << 94) +
      (src094[17] << 94) +
      (src094[18] << 94) +
      (src094[19] << 94) +
      (src094[20] << 94) +
      (src094[21] << 94) +
      (src094[22] << 94) +
      (src094[23] << 94) +
      (src094[24] << 94) +
      (src094[25] << 94) +
      (src094[26] << 94) +
      (src094[27] << 94) +
      (src094[28] << 94) +
      (src094[29] << 94) +
      (src094[30] << 94) +
      (src094[31] << 94) +
      (src094[32] << 94) +
      (src094[33] << 94) +
      (src094[34] << 94) +
      (src094[35] << 94) +
      (src094[36] << 94) +
      (src094[37] << 94) +
      (src094[38] << 94) +
      (src094[39] << 94) +
      (src094[40] << 94) +
      (src094[41] << 94) +
      (src094[42] << 94) +
      (src094[43] << 94) +
      (src094[44] << 94) +
      (src094[45] << 94) +
      (src094[46] << 94) +
      (src094[47] << 94) +
      (src094[48] << 94) +
      (src094[49] << 94) +
      (src094[50] << 94) +
      (src094[51] << 94) +
      (src094[52] << 94) +
      (src094[53] << 94) +
      (src094[54] << 94) +
      (src094[55] << 94) +
      (src094[56] << 94) +
      (src094[57] << 94) +
      (src094[58] << 94) +
      (src094[59] << 94) +
      (src094[60] << 94) +
      (src094[61] << 94) +
      (src094[62] << 94) +
      (src094[63] << 94) +
      (src094[64] << 94) +
      (src094[65] << 94) +
      (src094[66] << 94) +
      (src094[67] << 94) +
      (src094[68] << 94) +
      (src094[69] << 94) +
      (src094[70] << 94) +
      (src094[71] << 94) +
      (src094[72] << 94) +
      (src094[73] << 94) +
      (src094[74] << 94) +
      (src094[75] << 94) +
      (src094[76] << 94) +
      (src094[77] << 94) +
      (src094[78] << 94) +
      (src094[79] << 94) +
      (src094[80] << 94) +
      (src094[81] << 94) +
      (src094[82] << 94) +
      (src094[83] << 94) +
      (src094[84] << 94) +
      (src094[85] << 94) +
      (src094[86] << 94) +
      (src094[87] << 94) +
      (src094[88] << 94) +
      (src094[89] << 94) +
      (src094[90] << 94) +
      (src094[91] << 94) +
      (src094[92] << 94) +
      (src094[93] << 94) +
      (src094[94] << 94) +
      (src094[95] << 94) +
      (src094[96] << 94) +
      (src094[97] << 94) +
      (src094[98] << 94) +
      (src094[99] << 94) +
      (src094[100] << 94) +
      (src094[101] << 94) +
      (src094[102] << 94) +
      (src094[103] << 94) +
      (src094[104] << 94) +
      (src094[105] << 94) +
      (src094[106] << 94) +
      (src094[107] << 94) +
      (src094[108] << 94) +
      (src094[109] << 94) +
      (src094[110] << 94) +
      (src094[111] << 94) +
      (src094[112] << 94) +
      (src094[113] << 94) +
      (src094[114] << 94) +
      (src094[115] << 94) +
      (src094[116] << 94) +
      (src094[117] << 94) +
      (src094[118] << 94) +
      (src094[119] << 94) +
      (src094[120] << 94) +
      (src094[121] << 94) +
      (src094[122] << 94) +
      (src094[123] << 94) +
      (src094[124] << 94) +
      (src094[125] << 94) +
      (src094[126] << 94) +
      (src094[127] << 94) +
      (src095[0] << 95) +
      (src095[1] << 95) +
      (src095[2] << 95) +
      (src095[3] << 95) +
      (src095[4] << 95) +
      (src095[5] << 95) +
      (src095[6] << 95) +
      (src095[7] << 95) +
      (src095[8] << 95) +
      (src095[9] << 95) +
      (src095[10] << 95) +
      (src095[11] << 95) +
      (src095[12] << 95) +
      (src095[13] << 95) +
      (src095[14] << 95) +
      (src095[15] << 95) +
      (src095[16] << 95) +
      (src095[17] << 95) +
      (src095[18] << 95) +
      (src095[19] << 95) +
      (src095[20] << 95) +
      (src095[21] << 95) +
      (src095[22] << 95) +
      (src095[23] << 95) +
      (src095[24] << 95) +
      (src095[25] << 95) +
      (src095[26] << 95) +
      (src095[27] << 95) +
      (src095[28] << 95) +
      (src095[29] << 95) +
      (src095[30] << 95) +
      (src095[31] << 95) +
      (src095[32] << 95) +
      (src095[33] << 95) +
      (src095[34] << 95) +
      (src095[35] << 95) +
      (src095[36] << 95) +
      (src095[37] << 95) +
      (src095[38] << 95) +
      (src095[39] << 95) +
      (src095[40] << 95) +
      (src095[41] << 95) +
      (src095[42] << 95) +
      (src095[43] << 95) +
      (src095[44] << 95) +
      (src095[45] << 95) +
      (src095[46] << 95) +
      (src095[47] << 95) +
      (src095[48] << 95) +
      (src095[49] << 95) +
      (src095[50] << 95) +
      (src095[51] << 95) +
      (src095[52] << 95) +
      (src095[53] << 95) +
      (src095[54] << 95) +
      (src095[55] << 95) +
      (src095[56] << 95) +
      (src095[57] << 95) +
      (src095[58] << 95) +
      (src095[59] << 95) +
      (src095[60] << 95) +
      (src095[61] << 95) +
      (src095[62] << 95) +
      (src095[63] << 95) +
      (src095[64] << 95) +
      (src095[65] << 95) +
      (src095[66] << 95) +
      (src095[67] << 95) +
      (src095[68] << 95) +
      (src095[69] << 95) +
      (src095[70] << 95) +
      (src095[71] << 95) +
      (src095[72] << 95) +
      (src095[73] << 95) +
      (src095[74] << 95) +
      (src095[75] << 95) +
      (src095[76] << 95) +
      (src095[77] << 95) +
      (src095[78] << 95) +
      (src095[79] << 95) +
      (src095[80] << 95) +
      (src095[81] << 95) +
      (src095[82] << 95) +
      (src095[83] << 95) +
      (src095[84] << 95) +
      (src095[85] << 95) +
      (src095[86] << 95) +
      (src095[87] << 95) +
      (src095[88] << 95) +
      (src095[89] << 95) +
      (src095[90] << 95) +
      (src095[91] << 95) +
      (src095[92] << 95) +
      (src095[93] << 95) +
      (src095[94] << 95) +
      (src095[95] << 95) +
      (src095[96] << 95) +
      (src095[97] << 95) +
      (src095[98] << 95) +
      (src095[99] << 95) +
      (src095[100] << 95) +
      (src095[101] << 95) +
      (src095[102] << 95) +
      (src095[103] << 95) +
      (src095[104] << 95) +
      (src095[105] << 95) +
      (src095[106] << 95) +
      (src095[107] << 95) +
      (src095[108] << 95) +
      (src095[109] << 95) +
      (src095[110] << 95) +
      (src095[111] << 95) +
      (src095[112] << 95) +
      (src095[113] << 95) +
      (src095[114] << 95) +
      (src095[115] << 95) +
      (src095[116] << 95) +
      (src095[117] << 95) +
      (src095[118] << 95) +
      (src095[119] << 95) +
      (src095[120] << 95) +
      (src095[121] << 95) +
      (src095[122] << 95) +
      (src095[123] << 95) +
      (src095[124] << 95) +
      (src095[125] << 95) +
      (src095[126] << 95) +
      (src095[127] << 95) +
      (src096[0] << 96) +
      (src096[1] << 96) +
      (src096[2] << 96) +
      (src096[3] << 96) +
      (src096[4] << 96) +
      (src096[5] << 96) +
      (src096[6] << 96) +
      (src096[7] << 96) +
      (src096[8] << 96) +
      (src096[9] << 96) +
      (src096[10] << 96) +
      (src096[11] << 96) +
      (src096[12] << 96) +
      (src096[13] << 96) +
      (src096[14] << 96) +
      (src096[15] << 96) +
      (src096[16] << 96) +
      (src096[17] << 96) +
      (src096[18] << 96) +
      (src096[19] << 96) +
      (src096[20] << 96) +
      (src096[21] << 96) +
      (src096[22] << 96) +
      (src096[23] << 96) +
      (src096[24] << 96) +
      (src096[25] << 96) +
      (src096[26] << 96) +
      (src096[27] << 96) +
      (src096[28] << 96) +
      (src096[29] << 96) +
      (src096[30] << 96) +
      (src096[31] << 96) +
      (src096[32] << 96) +
      (src096[33] << 96) +
      (src096[34] << 96) +
      (src096[35] << 96) +
      (src096[36] << 96) +
      (src096[37] << 96) +
      (src096[38] << 96) +
      (src096[39] << 96) +
      (src096[40] << 96) +
      (src096[41] << 96) +
      (src096[42] << 96) +
      (src096[43] << 96) +
      (src096[44] << 96) +
      (src096[45] << 96) +
      (src096[46] << 96) +
      (src096[47] << 96) +
      (src096[48] << 96) +
      (src096[49] << 96) +
      (src096[50] << 96) +
      (src096[51] << 96) +
      (src096[52] << 96) +
      (src096[53] << 96) +
      (src096[54] << 96) +
      (src096[55] << 96) +
      (src096[56] << 96) +
      (src096[57] << 96) +
      (src096[58] << 96) +
      (src096[59] << 96) +
      (src096[60] << 96) +
      (src096[61] << 96) +
      (src096[62] << 96) +
      (src096[63] << 96) +
      (src096[64] << 96) +
      (src096[65] << 96) +
      (src096[66] << 96) +
      (src096[67] << 96) +
      (src096[68] << 96) +
      (src096[69] << 96) +
      (src096[70] << 96) +
      (src096[71] << 96) +
      (src096[72] << 96) +
      (src096[73] << 96) +
      (src096[74] << 96) +
      (src096[75] << 96) +
      (src096[76] << 96) +
      (src096[77] << 96) +
      (src096[78] << 96) +
      (src096[79] << 96) +
      (src096[80] << 96) +
      (src096[81] << 96) +
      (src096[82] << 96) +
      (src096[83] << 96) +
      (src096[84] << 96) +
      (src096[85] << 96) +
      (src096[86] << 96) +
      (src096[87] << 96) +
      (src096[88] << 96) +
      (src096[89] << 96) +
      (src096[90] << 96) +
      (src096[91] << 96) +
      (src096[92] << 96) +
      (src096[93] << 96) +
      (src096[94] << 96) +
      (src096[95] << 96) +
      (src096[96] << 96) +
      (src096[97] << 96) +
      (src096[98] << 96) +
      (src096[99] << 96) +
      (src096[100] << 96) +
      (src096[101] << 96) +
      (src096[102] << 96) +
      (src096[103] << 96) +
      (src096[104] << 96) +
      (src096[105] << 96) +
      (src096[106] << 96) +
      (src096[107] << 96) +
      (src096[108] << 96) +
      (src096[109] << 96) +
      (src096[110] << 96) +
      (src096[111] << 96) +
      (src096[112] << 96) +
      (src096[113] << 96) +
      (src096[114] << 96) +
      (src096[115] << 96) +
      (src096[116] << 96) +
      (src096[117] << 96) +
      (src096[118] << 96) +
      (src096[119] << 96) +
      (src096[120] << 96) +
      (src096[121] << 96) +
      (src096[122] << 96) +
      (src096[123] << 96) +
      (src096[124] << 96) +
      (src096[125] << 96) +
      (src096[126] << 96) +
      (src096[127] << 96) +
      (src097[0] << 97) +
      (src097[1] << 97) +
      (src097[2] << 97) +
      (src097[3] << 97) +
      (src097[4] << 97) +
      (src097[5] << 97) +
      (src097[6] << 97) +
      (src097[7] << 97) +
      (src097[8] << 97) +
      (src097[9] << 97) +
      (src097[10] << 97) +
      (src097[11] << 97) +
      (src097[12] << 97) +
      (src097[13] << 97) +
      (src097[14] << 97) +
      (src097[15] << 97) +
      (src097[16] << 97) +
      (src097[17] << 97) +
      (src097[18] << 97) +
      (src097[19] << 97) +
      (src097[20] << 97) +
      (src097[21] << 97) +
      (src097[22] << 97) +
      (src097[23] << 97) +
      (src097[24] << 97) +
      (src097[25] << 97) +
      (src097[26] << 97) +
      (src097[27] << 97) +
      (src097[28] << 97) +
      (src097[29] << 97) +
      (src097[30] << 97) +
      (src097[31] << 97) +
      (src097[32] << 97) +
      (src097[33] << 97) +
      (src097[34] << 97) +
      (src097[35] << 97) +
      (src097[36] << 97) +
      (src097[37] << 97) +
      (src097[38] << 97) +
      (src097[39] << 97) +
      (src097[40] << 97) +
      (src097[41] << 97) +
      (src097[42] << 97) +
      (src097[43] << 97) +
      (src097[44] << 97) +
      (src097[45] << 97) +
      (src097[46] << 97) +
      (src097[47] << 97) +
      (src097[48] << 97) +
      (src097[49] << 97) +
      (src097[50] << 97) +
      (src097[51] << 97) +
      (src097[52] << 97) +
      (src097[53] << 97) +
      (src097[54] << 97) +
      (src097[55] << 97) +
      (src097[56] << 97) +
      (src097[57] << 97) +
      (src097[58] << 97) +
      (src097[59] << 97) +
      (src097[60] << 97) +
      (src097[61] << 97) +
      (src097[62] << 97) +
      (src097[63] << 97) +
      (src097[64] << 97) +
      (src097[65] << 97) +
      (src097[66] << 97) +
      (src097[67] << 97) +
      (src097[68] << 97) +
      (src097[69] << 97) +
      (src097[70] << 97) +
      (src097[71] << 97) +
      (src097[72] << 97) +
      (src097[73] << 97) +
      (src097[74] << 97) +
      (src097[75] << 97) +
      (src097[76] << 97) +
      (src097[77] << 97) +
      (src097[78] << 97) +
      (src097[79] << 97) +
      (src097[80] << 97) +
      (src097[81] << 97) +
      (src097[82] << 97) +
      (src097[83] << 97) +
      (src097[84] << 97) +
      (src097[85] << 97) +
      (src097[86] << 97) +
      (src097[87] << 97) +
      (src097[88] << 97) +
      (src097[89] << 97) +
      (src097[90] << 97) +
      (src097[91] << 97) +
      (src097[92] << 97) +
      (src097[93] << 97) +
      (src097[94] << 97) +
      (src097[95] << 97) +
      (src097[96] << 97) +
      (src097[97] << 97) +
      (src097[98] << 97) +
      (src097[99] << 97) +
      (src097[100] << 97) +
      (src097[101] << 97) +
      (src097[102] << 97) +
      (src097[103] << 97) +
      (src097[104] << 97) +
      (src097[105] << 97) +
      (src097[106] << 97) +
      (src097[107] << 97) +
      (src097[108] << 97) +
      (src097[109] << 97) +
      (src097[110] << 97) +
      (src097[111] << 97) +
      (src097[112] << 97) +
      (src097[113] << 97) +
      (src097[114] << 97) +
      (src097[115] << 97) +
      (src097[116] << 97) +
      (src097[117] << 97) +
      (src097[118] << 97) +
      (src097[119] << 97) +
      (src097[120] << 97) +
      (src097[121] << 97) +
      (src097[122] << 97) +
      (src097[123] << 97) +
      (src097[124] << 97) +
      (src097[125] << 97) +
      (src097[126] << 97) +
      (src097[127] << 97) +
      (src098[0] << 98) +
      (src098[1] << 98) +
      (src098[2] << 98) +
      (src098[3] << 98) +
      (src098[4] << 98) +
      (src098[5] << 98) +
      (src098[6] << 98) +
      (src098[7] << 98) +
      (src098[8] << 98) +
      (src098[9] << 98) +
      (src098[10] << 98) +
      (src098[11] << 98) +
      (src098[12] << 98) +
      (src098[13] << 98) +
      (src098[14] << 98) +
      (src098[15] << 98) +
      (src098[16] << 98) +
      (src098[17] << 98) +
      (src098[18] << 98) +
      (src098[19] << 98) +
      (src098[20] << 98) +
      (src098[21] << 98) +
      (src098[22] << 98) +
      (src098[23] << 98) +
      (src098[24] << 98) +
      (src098[25] << 98) +
      (src098[26] << 98) +
      (src098[27] << 98) +
      (src098[28] << 98) +
      (src098[29] << 98) +
      (src098[30] << 98) +
      (src098[31] << 98) +
      (src098[32] << 98) +
      (src098[33] << 98) +
      (src098[34] << 98) +
      (src098[35] << 98) +
      (src098[36] << 98) +
      (src098[37] << 98) +
      (src098[38] << 98) +
      (src098[39] << 98) +
      (src098[40] << 98) +
      (src098[41] << 98) +
      (src098[42] << 98) +
      (src098[43] << 98) +
      (src098[44] << 98) +
      (src098[45] << 98) +
      (src098[46] << 98) +
      (src098[47] << 98) +
      (src098[48] << 98) +
      (src098[49] << 98) +
      (src098[50] << 98) +
      (src098[51] << 98) +
      (src098[52] << 98) +
      (src098[53] << 98) +
      (src098[54] << 98) +
      (src098[55] << 98) +
      (src098[56] << 98) +
      (src098[57] << 98) +
      (src098[58] << 98) +
      (src098[59] << 98) +
      (src098[60] << 98) +
      (src098[61] << 98) +
      (src098[62] << 98) +
      (src098[63] << 98) +
      (src098[64] << 98) +
      (src098[65] << 98) +
      (src098[66] << 98) +
      (src098[67] << 98) +
      (src098[68] << 98) +
      (src098[69] << 98) +
      (src098[70] << 98) +
      (src098[71] << 98) +
      (src098[72] << 98) +
      (src098[73] << 98) +
      (src098[74] << 98) +
      (src098[75] << 98) +
      (src098[76] << 98) +
      (src098[77] << 98) +
      (src098[78] << 98) +
      (src098[79] << 98) +
      (src098[80] << 98) +
      (src098[81] << 98) +
      (src098[82] << 98) +
      (src098[83] << 98) +
      (src098[84] << 98) +
      (src098[85] << 98) +
      (src098[86] << 98) +
      (src098[87] << 98) +
      (src098[88] << 98) +
      (src098[89] << 98) +
      (src098[90] << 98) +
      (src098[91] << 98) +
      (src098[92] << 98) +
      (src098[93] << 98) +
      (src098[94] << 98) +
      (src098[95] << 98) +
      (src098[96] << 98) +
      (src098[97] << 98) +
      (src098[98] << 98) +
      (src098[99] << 98) +
      (src098[100] << 98) +
      (src098[101] << 98) +
      (src098[102] << 98) +
      (src098[103] << 98) +
      (src098[104] << 98) +
      (src098[105] << 98) +
      (src098[106] << 98) +
      (src098[107] << 98) +
      (src098[108] << 98) +
      (src098[109] << 98) +
      (src098[110] << 98) +
      (src098[111] << 98) +
      (src098[112] << 98) +
      (src098[113] << 98) +
      (src098[114] << 98) +
      (src098[115] << 98) +
      (src098[116] << 98) +
      (src098[117] << 98) +
      (src098[118] << 98) +
      (src098[119] << 98) +
      (src098[120] << 98) +
      (src098[121] << 98) +
      (src098[122] << 98) +
      (src098[123] << 98) +
      (src098[124] << 98) +
      (src098[125] << 98) +
      (src098[126] << 98) +
      (src098[127] << 98) +
      (src099[0] << 99) +
      (src099[1] << 99) +
      (src099[2] << 99) +
      (src099[3] << 99) +
      (src099[4] << 99) +
      (src099[5] << 99) +
      (src099[6] << 99) +
      (src099[7] << 99) +
      (src099[8] << 99) +
      (src099[9] << 99) +
      (src099[10] << 99) +
      (src099[11] << 99) +
      (src099[12] << 99) +
      (src099[13] << 99) +
      (src099[14] << 99) +
      (src099[15] << 99) +
      (src099[16] << 99) +
      (src099[17] << 99) +
      (src099[18] << 99) +
      (src099[19] << 99) +
      (src099[20] << 99) +
      (src099[21] << 99) +
      (src099[22] << 99) +
      (src099[23] << 99) +
      (src099[24] << 99) +
      (src099[25] << 99) +
      (src099[26] << 99) +
      (src099[27] << 99) +
      (src099[28] << 99) +
      (src099[29] << 99) +
      (src099[30] << 99) +
      (src099[31] << 99) +
      (src099[32] << 99) +
      (src099[33] << 99) +
      (src099[34] << 99) +
      (src099[35] << 99) +
      (src099[36] << 99) +
      (src099[37] << 99) +
      (src099[38] << 99) +
      (src099[39] << 99) +
      (src099[40] << 99) +
      (src099[41] << 99) +
      (src099[42] << 99) +
      (src099[43] << 99) +
      (src099[44] << 99) +
      (src099[45] << 99) +
      (src099[46] << 99) +
      (src099[47] << 99) +
      (src099[48] << 99) +
      (src099[49] << 99) +
      (src099[50] << 99) +
      (src099[51] << 99) +
      (src099[52] << 99) +
      (src099[53] << 99) +
      (src099[54] << 99) +
      (src099[55] << 99) +
      (src099[56] << 99) +
      (src099[57] << 99) +
      (src099[58] << 99) +
      (src099[59] << 99) +
      (src099[60] << 99) +
      (src099[61] << 99) +
      (src099[62] << 99) +
      (src099[63] << 99) +
      (src099[64] << 99) +
      (src099[65] << 99) +
      (src099[66] << 99) +
      (src099[67] << 99) +
      (src099[68] << 99) +
      (src099[69] << 99) +
      (src099[70] << 99) +
      (src099[71] << 99) +
      (src099[72] << 99) +
      (src099[73] << 99) +
      (src099[74] << 99) +
      (src099[75] << 99) +
      (src099[76] << 99) +
      (src099[77] << 99) +
      (src099[78] << 99) +
      (src099[79] << 99) +
      (src099[80] << 99) +
      (src099[81] << 99) +
      (src099[82] << 99) +
      (src099[83] << 99) +
      (src099[84] << 99) +
      (src099[85] << 99) +
      (src099[86] << 99) +
      (src099[87] << 99) +
      (src099[88] << 99) +
      (src099[89] << 99) +
      (src099[90] << 99) +
      (src099[91] << 99) +
      (src099[92] << 99) +
      (src099[93] << 99) +
      (src099[94] << 99) +
      (src099[95] << 99) +
      (src099[96] << 99) +
      (src099[97] << 99) +
      (src099[98] << 99) +
      (src099[99] << 99) +
      (src099[100] << 99) +
      (src099[101] << 99) +
      (src099[102] << 99) +
      (src099[103] << 99) +
      (src099[104] << 99) +
      (src099[105] << 99) +
      (src099[106] << 99) +
      (src099[107] << 99) +
      (src099[108] << 99) +
      (src099[109] << 99) +
      (src099[110] << 99) +
      (src099[111] << 99) +
      (src099[112] << 99) +
      (src099[113] << 99) +
      (src099[114] << 99) +
      (src099[115] << 99) +
      (src099[116] << 99) +
      (src099[117] << 99) +
      (src099[118] << 99) +
      (src099[119] << 99) +
      (src099[120] << 99) +
      (src099[121] << 99) +
      (src099[122] << 99) +
      (src099[123] << 99) +
      (src099[124] << 99) +
      (src099[125] << 99) +
      (src099[126] << 99) +
      (src099[127] << 99) +
      (src100[0] << 100) +
      (src100[1] << 100) +
      (src100[2] << 100) +
      (src100[3] << 100) +
      (src100[4] << 100) +
      (src100[5] << 100) +
      (src100[6] << 100) +
      (src100[7] << 100) +
      (src100[8] << 100) +
      (src100[9] << 100) +
      (src100[10] << 100) +
      (src100[11] << 100) +
      (src100[12] << 100) +
      (src100[13] << 100) +
      (src100[14] << 100) +
      (src100[15] << 100) +
      (src100[16] << 100) +
      (src100[17] << 100) +
      (src100[18] << 100) +
      (src100[19] << 100) +
      (src100[20] << 100) +
      (src100[21] << 100) +
      (src100[22] << 100) +
      (src100[23] << 100) +
      (src100[24] << 100) +
      (src100[25] << 100) +
      (src100[26] << 100) +
      (src100[27] << 100) +
      (src100[28] << 100) +
      (src100[29] << 100) +
      (src100[30] << 100) +
      (src100[31] << 100) +
      (src100[32] << 100) +
      (src100[33] << 100) +
      (src100[34] << 100) +
      (src100[35] << 100) +
      (src100[36] << 100) +
      (src100[37] << 100) +
      (src100[38] << 100) +
      (src100[39] << 100) +
      (src100[40] << 100) +
      (src100[41] << 100) +
      (src100[42] << 100) +
      (src100[43] << 100) +
      (src100[44] << 100) +
      (src100[45] << 100) +
      (src100[46] << 100) +
      (src100[47] << 100) +
      (src100[48] << 100) +
      (src100[49] << 100) +
      (src100[50] << 100) +
      (src100[51] << 100) +
      (src100[52] << 100) +
      (src100[53] << 100) +
      (src100[54] << 100) +
      (src100[55] << 100) +
      (src100[56] << 100) +
      (src100[57] << 100) +
      (src100[58] << 100) +
      (src100[59] << 100) +
      (src100[60] << 100) +
      (src100[61] << 100) +
      (src100[62] << 100) +
      (src100[63] << 100) +
      (src100[64] << 100) +
      (src100[65] << 100) +
      (src100[66] << 100) +
      (src100[67] << 100) +
      (src100[68] << 100) +
      (src100[69] << 100) +
      (src100[70] << 100) +
      (src100[71] << 100) +
      (src100[72] << 100) +
      (src100[73] << 100) +
      (src100[74] << 100) +
      (src100[75] << 100) +
      (src100[76] << 100) +
      (src100[77] << 100) +
      (src100[78] << 100) +
      (src100[79] << 100) +
      (src100[80] << 100) +
      (src100[81] << 100) +
      (src100[82] << 100) +
      (src100[83] << 100) +
      (src100[84] << 100) +
      (src100[85] << 100) +
      (src100[86] << 100) +
      (src100[87] << 100) +
      (src100[88] << 100) +
      (src100[89] << 100) +
      (src100[90] << 100) +
      (src100[91] << 100) +
      (src100[92] << 100) +
      (src100[93] << 100) +
      (src100[94] << 100) +
      (src100[95] << 100) +
      (src100[96] << 100) +
      (src100[97] << 100) +
      (src100[98] << 100) +
      (src100[99] << 100) +
      (src100[100] << 100) +
      (src100[101] << 100) +
      (src100[102] << 100) +
      (src100[103] << 100) +
      (src100[104] << 100) +
      (src100[105] << 100) +
      (src100[106] << 100) +
      (src100[107] << 100) +
      (src100[108] << 100) +
      (src100[109] << 100) +
      (src100[110] << 100) +
      (src100[111] << 100) +
      (src100[112] << 100) +
      (src100[113] << 100) +
      (src100[114] << 100) +
      (src100[115] << 100) +
      (src100[116] << 100) +
      (src100[117] << 100) +
      (src100[118] << 100) +
      (src100[119] << 100) +
      (src100[120] << 100) +
      (src100[121] << 100) +
      (src100[122] << 100) +
      (src100[123] << 100) +
      (src100[124] << 100) +
      (src100[125] << 100) +
      (src100[126] << 100) +
      (src100[127] << 100) +
      (src101[0] << 101) +
      (src101[1] << 101) +
      (src101[2] << 101) +
      (src101[3] << 101) +
      (src101[4] << 101) +
      (src101[5] << 101) +
      (src101[6] << 101) +
      (src101[7] << 101) +
      (src101[8] << 101) +
      (src101[9] << 101) +
      (src101[10] << 101) +
      (src101[11] << 101) +
      (src101[12] << 101) +
      (src101[13] << 101) +
      (src101[14] << 101) +
      (src101[15] << 101) +
      (src101[16] << 101) +
      (src101[17] << 101) +
      (src101[18] << 101) +
      (src101[19] << 101) +
      (src101[20] << 101) +
      (src101[21] << 101) +
      (src101[22] << 101) +
      (src101[23] << 101) +
      (src101[24] << 101) +
      (src101[25] << 101) +
      (src101[26] << 101) +
      (src101[27] << 101) +
      (src101[28] << 101) +
      (src101[29] << 101) +
      (src101[30] << 101) +
      (src101[31] << 101) +
      (src101[32] << 101) +
      (src101[33] << 101) +
      (src101[34] << 101) +
      (src101[35] << 101) +
      (src101[36] << 101) +
      (src101[37] << 101) +
      (src101[38] << 101) +
      (src101[39] << 101) +
      (src101[40] << 101) +
      (src101[41] << 101) +
      (src101[42] << 101) +
      (src101[43] << 101) +
      (src101[44] << 101) +
      (src101[45] << 101) +
      (src101[46] << 101) +
      (src101[47] << 101) +
      (src101[48] << 101) +
      (src101[49] << 101) +
      (src101[50] << 101) +
      (src101[51] << 101) +
      (src101[52] << 101) +
      (src101[53] << 101) +
      (src101[54] << 101) +
      (src101[55] << 101) +
      (src101[56] << 101) +
      (src101[57] << 101) +
      (src101[58] << 101) +
      (src101[59] << 101) +
      (src101[60] << 101) +
      (src101[61] << 101) +
      (src101[62] << 101) +
      (src101[63] << 101) +
      (src101[64] << 101) +
      (src101[65] << 101) +
      (src101[66] << 101) +
      (src101[67] << 101) +
      (src101[68] << 101) +
      (src101[69] << 101) +
      (src101[70] << 101) +
      (src101[71] << 101) +
      (src101[72] << 101) +
      (src101[73] << 101) +
      (src101[74] << 101) +
      (src101[75] << 101) +
      (src101[76] << 101) +
      (src101[77] << 101) +
      (src101[78] << 101) +
      (src101[79] << 101) +
      (src101[80] << 101) +
      (src101[81] << 101) +
      (src101[82] << 101) +
      (src101[83] << 101) +
      (src101[84] << 101) +
      (src101[85] << 101) +
      (src101[86] << 101) +
      (src101[87] << 101) +
      (src101[88] << 101) +
      (src101[89] << 101) +
      (src101[90] << 101) +
      (src101[91] << 101) +
      (src101[92] << 101) +
      (src101[93] << 101) +
      (src101[94] << 101) +
      (src101[95] << 101) +
      (src101[96] << 101) +
      (src101[97] << 101) +
      (src101[98] << 101) +
      (src101[99] << 101) +
      (src101[100] << 101) +
      (src101[101] << 101) +
      (src101[102] << 101) +
      (src101[103] << 101) +
      (src101[104] << 101) +
      (src101[105] << 101) +
      (src101[106] << 101) +
      (src101[107] << 101) +
      (src101[108] << 101) +
      (src101[109] << 101) +
      (src101[110] << 101) +
      (src101[111] << 101) +
      (src101[112] << 101) +
      (src101[113] << 101) +
      (src101[114] << 101) +
      (src101[115] << 101) +
      (src101[116] << 101) +
      (src101[117] << 101) +
      (src101[118] << 101) +
      (src101[119] << 101) +
      (src101[120] << 101) +
      (src101[121] << 101) +
      (src101[122] << 101) +
      (src101[123] << 101) +
      (src101[124] << 101) +
      (src101[125] << 101) +
      (src101[126] << 101) +
      (src101[127] << 101) +
      (src102[0] << 102) +
      (src102[1] << 102) +
      (src102[2] << 102) +
      (src102[3] << 102) +
      (src102[4] << 102) +
      (src102[5] << 102) +
      (src102[6] << 102) +
      (src102[7] << 102) +
      (src102[8] << 102) +
      (src102[9] << 102) +
      (src102[10] << 102) +
      (src102[11] << 102) +
      (src102[12] << 102) +
      (src102[13] << 102) +
      (src102[14] << 102) +
      (src102[15] << 102) +
      (src102[16] << 102) +
      (src102[17] << 102) +
      (src102[18] << 102) +
      (src102[19] << 102) +
      (src102[20] << 102) +
      (src102[21] << 102) +
      (src102[22] << 102) +
      (src102[23] << 102) +
      (src102[24] << 102) +
      (src102[25] << 102) +
      (src102[26] << 102) +
      (src102[27] << 102) +
      (src102[28] << 102) +
      (src102[29] << 102) +
      (src102[30] << 102) +
      (src102[31] << 102) +
      (src102[32] << 102) +
      (src102[33] << 102) +
      (src102[34] << 102) +
      (src102[35] << 102) +
      (src102[36] << 102) +
      (src102[37] << 102) +
      (src102[38] << 102) +
      (src102[39] << 102) +
      (src102[40] << 102) +
      (src102[41] << 102) +
      (src102[42] << 102) +
      (src102[43] << 102) +
      (src102[44] << 102) +
      (src102[45] << 102) +
      (src102[46] << 102) +
      (src102[47] << 102) +
      (src102[48] << 102) +
      (src102[49] << 102) +
      (src102[50] << 102) +
      (src102[51] << 102) +
      (src102[52] << 102) +
      (src102[53] << 102) +
      (src102[54] << 102) +
      (src102[55] << 102) +
      (src102[56] << 102) +
      (src102[57] << 102) +
      (src102[58] << 102) +
      (src102[59] << 102) +
      (src102[60] << 102) +
      (src102[61] << 102) +
      (src102[62] << 102) +
      (src102[63] << 102) +
      (src102[64] << 102) +
      (src102[65] << 102) +
      (src102[66] << 102) +
      (src102[67] << 102) +
      (src102[68] << 102) +
      (src102[69] << 102) +
      (src102[70] << 102) +
      (src102[71] << 102) +
      (src102[72] << 102) +
      (src102[73] << 102) +
      (src102[74] << 102) +
      (src102[75] << 102) +
      (src102[76] << 102) +
      (src102[77] << 102) +
      (src102[78] << 102) +
      (src102[79] << 102) +
      (src102[80] << 102) +
      (src102[81] << 102) +
      (src102[82] << 102) +
      (src102[83] << 102) +
      (src102[84] << 102) +
      (src102[85] << 102) +
      (src102[86] << 102) +
      (src102[87] << 102) +
      (src102[88] << 102) +
      (src102[89] << 102) +
      (src102[90] << 102) +
      (src102[91] << 102) +
      (src102[92] << 102) +
      (src102[93] << 102) +
      (src102[94] << 102) +
      (src102[95] << 102) +
      (src102[96] << 102) +
      (src102[97] << 102) +
      (src102[98] << 102) +
      (src102[99] << 102) +
      (src102[100] << 102) +
      (src102[101] << 102) +
      (src102[102] << 102) +
      (src102[103] << 102) +
      (src102[104] << 102) +
      (src102[105] << 102) +
      (src102[106] << 102) +
      (src102[107] << 102) +
      (src102[108] << 102) +
      (src102[109] << 102) +
      (src102[110] << 102) +
      (src102[111] << 102) +
      (src102[112] << 102) +
      (src102[113] << 102) +
      (src102[114] << 102) +
      (src102[115] << 102) +
      (src102[116] << 102) +
      (src102[117] << 102) +
      (src102[118] << 102) +
      (src102[119] << 102) +
      (src102[120] << 102) +
      (src102[121] << 102) +
      (src102[122] << 102) +
      (src102[123] << 102) +
      (src102[124] << 102) +
      (src102[125] << 102) +
      (src102[126] << 102) +
      (src102[127] << 102) +
      (src103[0] << 103) +
      (src103[1] << 103) +
      (src103[2] << 103) +
      (src103[3] << 103) +
      (src103[4] << 103) +
      (src103[5] << 103) +
      (src103[6] << 103) +
      (src103[7] << 103) +
      (src103[8] << 103) +
      (src103[9] << 103) +
      (src103[10] << 103) +
      (src103[11] << 103) +
      (src103[12] << 103) +
      (src103[13] << 103) +
      (src103[14] << 103) +
      (src103[15] << 103) +
      (src103[16] << 103) +
      (src103[17] << 103) +
      (src103[18] << 103) +
      (src103[19] << 103) +
      (src103[20] << 103) +
      (src103[21] << 103) +
      (src103[22] << 103) +
      (src103[23] << 103) +
      (src103[24] << 103) +
      (src103[25] << 103) +
      (src103[26] << 103) +
      (src103[27] << 103) +
      (src103[28] << 103) +
      (src103[29] << 103) +
      (src103[30] << 103) +
      (src103[31] << 103) +
      (src103[32] << 103) +
      (src103[33] << 103) +
      (src103[34] << 103) +
      (src103[35] << 103) +
      (src103[36] << 103) +
      (src103[37] << 103) +
      (src103[38] << 103) +
      (src103[39] << 103) +
      (src103[40] << 103) +
      (src103[41] << 103) +
      (src103[42] << 103) +
      (src103[43] << 103) +
      (src103[44] << 103) +
      (src103[45] << 103) +
      (src103[46] << 103) +
      (src103[47] << 103) +
      (src103[48] << 103) +
      (src103[49] << 103) +
      (src103[50] << 103) +
      (src103[51] << 103) +
      (src103[52] << 103) +
      (src103[53] << 103) +
      (src103[54] << 103) +
      (src103[55] << 103) +
      (src103[56] << 103) +
      (src103[57] << 103) +
      (src103[58] << 103) +
      (src103[59] << 103) +
      (src103[60] << 103) +
      (src103[61] << 103) +
      (src103[62] << 103) +
      (src103[63] << 103) +
      (src103[64] << 103) +
      (src103[65] << 103) +
      (src103[66] << 103) +
      (src103[67] << 103) +
      (src103[68] << 103) +
      (src103[69] << 103) +
      (src103[70] << 103) +
      (src103[71] << 103) +
      (src103[72] << 103) +
      (src103[73] << 103) +
      (src103[74] << 103) +
      (src103[75] << 103) +
      (src103[76] << 103) +
      (src103[77] << 103) +
      (src103[78] << 103) +
      (src103[79] << 103) +
      (src103[80] << 103) +
      (src103[81] << 103) +
      (src103[82] << 103) +
      (src103[83] << 103) +
      (src103[84] << 103) +
      (src103[85] << 103) +
      (src103[86] << 103) +
      (src103[87] << 103) +
      (src103[88] << 103) +
      (src103[89] << 103) +
      (src103[90] << 103) +
      (src103[91] << 103) +
      (src103[92] << 103) +
      (src103[93] << 103) +
      (src103[94] << 103) +
      (src103[95] << 103) +
      (src103[96] << 103) +
      (src103[97] << 103) +
      (src103[98] << 103) +
      (src103[99] << 103) +
      (src103[100] << 103) +
      (src103[101] << 103) +
      (src103[102] << 103) +
      (src103[103] << 103) +
      (src103[104] << 103) +
      (src103[105] << 103) +
      (src103[106] << 103) +
      (src103[107] << 103) +
      (src103[108] << 103) +
      (src103[109] << 103) +
      (src103[110] << 103) +
      (src103[111] << 103) +
      (src103[112] << 103) +
      (src103[113] << 103) +
      (src103[114] << 103) +
      (src103[115] << 103) +
      (src103[116] << 103) +
      (src103[117] << 103) +
      (src103[118] << 103) +
      (src103[119] << 103) +
      (src103[120] << 103) +
      (src103[121] << 103) +
      (src103[122] << 103) +
      (src103[123] << 103) +
      (src103[124] << 103) +
      (src103[125] << 103) +
      (src103[126] << 103) +
      (src103[127] << 103) +
      (src104[0] << 104) +
      (src104[1] << 104) +
      (src104[2] << 104) +
      (src104[3] << 104) +
      (src104[4] << 104) +
      (src104[5] << 104) +
      (src104[6] << 104) +
      (src104[7] << 104) +
      (src104[8] << 104) +
      (src104[9] << 104) +
      (src104[10] << 104) +
      (src104[11] << 104) +
      (src104[12] << 104) +
      (src104[13] << 104) +
      (src104[14] << 104) +
      (src104[15] << 104) +
      (src104[16] << 104) +
      (src104[17] << 104) +
      (src104[18] << 104) +
      (src104[19] << 104) +
      (src104[20] << 104) +
      (src104[21] << 104) +
      (src104[22] << 104) +
      (src104[23] << 104) +
      (src104[24] << 104) +
      (src104[25] << 104) +
      (src104[26] << 104) +
      (src104[27] << 104) +
      (src104[28] << 104) +
      (src104[29] << 104) +
      (src104[30] << 104) +
      (src104[31] << 104) +
      (src104[32] << 104) +
      (src104[33] << 104) +
      (src104[34] << 104) +
      (src104[35] << 104) +
      (src104[36] << 104) +
      (src104[37] << 104) +
      (src104[38] << 104) +
      (src104[39] << 104) +
      (src104[40] << 104) +
      (src104[41] << 104) +
      (src104[42] << 104) +
      (src104[43] << 104) +
      (src104[44] << 104) +
      (src104[45] << 104) +
      (src104[46] << 104) +
      (src104[47] << 104) +
      (src104[48] << 104) +
      (src104[49] << 104) +
      (src104[50] << 104) +
      (src104[51] << 104) +
      (src104[52] << 104) +
      (src104[53] << 104) +
      (src104[54] << 104) +
      (src104[55] << 104) +
      (src104[56] << 104) +
      (src104[57] << 104) +
      (src104[58] << 104) +
      (src104[59] << 104) +
      (src104[60] << 104) +
      (src104[61] << 104) +
      (src104[62] << 104) +
      (src104[63] << 104) +
      (src104[64] << 104) +
      (src104[65] << 104) +
      (src104[66] << 104) +
      (src104[67] << 104) +
      (src104[68] << 104) +
      (src104[69] << 104) +
      (src104[70] << 104) +
      (src104[71] << 104) +
      (src104[72] << 104) +
      (src104[73] << 104) +
      (src104[74] << 104) +
      (src104[75] << 104) +
      (src104[76] << 104) +
      (src104[77] << 104) +
      (src104[78] << 104) +
      (src104[79] << 104) +
      (src104[80] << 104) +
      (src104[81] << 104) +
      (src104[82] << 104) +
      (src104[83] << 104) +
      (src104[84] << 104) +
      (src104[85] << 104) +
      (src104[86] << 104) +
      (src104[87] << 104) +
      (src104[88] << 104) +
      (src104[89] << 104) +
      (src104[90] << 104) +
      (src104[91] << 104) +
      (src104[92] << 104) +
      (src104[93] << 104) +
      (src104[94] << 104) +
      (src104[95] << 104) +
      (src104[96] << 104) +
      (src104[97] << 104) +
      (src104[98] << 104) +
      (src104[99] << 104) +
      (src104[100] << 104) +
      (src104[101] << 104) +
      (src104[102] << 104) +
      (src104[103] << 104) +
      (src104[104] << 104) +
      (src104[105] << 104) +
      (src104[106] << 104) +
      (src104[107] << 104) +
      (src104[108] << 104) +
      (src104[109] << 104) +
      (src104[110] << 104) +
      (src104[111] << 104) +
      (src104[112] << 104) +
      (src104[113] << 104) +
      (src104[114] << 104) +
      (src104[115] << 104) +
      (src104[116] << 104) +
      (src104[117] << 104) +
      (src104[118] << 104) +
      (src104[119] << 104) +
      (src104[120] << 104) +
      (src104[121] << 104) +
      (src104[122] << 104) +
      (src104[123] << 104) +
      (src104[124] << 104) +
      (src104[125] << 104) +
      (src104[126] << 104) +
      (src104[127] << 104) +
      (src105[0] << 105) +
      (src105[1] << 105) +
      (src105[2] << 105) +
      (src105[3] << 105) +
      (src105[4] << 105) +
      (src105[5] << 105) +
      (src105[6] << 105) +
      (src105[7] << 105) +
      (src105[8] << 105) +
      (src105[9] << 105) +
      (src105[10] << 105) +
      (src105[11] << 105) +
      (src105[12] << 105) +
      (src105[13] << 105) +
      (src105[14] << 105) +
      (src105[15] << 105) +
      (src105[16] << 105) +
      (src105[17] << 105) +
      (src105[18] << 105) +
      (src105[19] << 105) +
      (src105[20] << 105) +
      (src105[21] << 105) +
      (src105[22] << 105) +
      (src105[23] << 105) +
      (src105[24] << 105) +
      (src105[25] << 105) +
      (src105[26] << 105) +
      (src105[27] << 105) +
      (src105[28] << 105) +
      (src105[29] << 105) +
      (src105[30] << 105) +
      (src105[31] << 105) +
      (src105[32] << 105) +
      (src105[33] << 105) +
      (src105[34] << 105) +
      (src105[35] << 105) +
      (src105[36] << 105) +
      (src105[37] << 105) +
      (src105[38] << 105) +
      (src105[39] << 105) +
      (src105[40] << 105) +
      (src105[41] << 105) +
      (src105[42] << 105) +
      (src105[43] << 105) +
      (src105[44] << 105) +
      (src105[45] << 105) +
      (src105[46] << 105) +
      (src105[47] << 105) +
      (src105[48] << 105) +
      (src105[49] << 105) +
      (src105[50] << 105) +
      (src105[51] << 105) +
      (src105[52] << 105) +
      (src105[53] << 105) +
      (src105[54] << 105) +
      (src105[55] << 105) +
      (src105[56] << 105) +
      (src105[57] << 105) +
      (src105[58] << 105) +
      (src105[59] << 105) +
      (src105[60] << 105) +
      (src105[61] << 105) +
      (src105[62] << 105) +
      (src105[63] << 105) +
      (src105[64] << 105) +
      (src105[65] << 105) +
      (src105[66] << 105) +
      (src105[67] << 105) +
      (src105[68] << 105) +
      (src105[69] << 105) +
      (src105[70] << 105) +
      (src105[71] << 105) +
      (src105[72] << 105) +
      (src105[73] << 105) +
      (src105[74] << 105) +
      (src105[75] << 105) +
      (src105[76] << 105) +
      (src105[77] << 105) +
      (src105[78] << 105) +
      (src105[79] << 105) +
      (src105[80] << 105) +
      (src105[81] << 105) +
      (src105[82] << 105) +
      (src105[83] << 105) +
      (src105[84] << 105) +
      (src105[85] << 105) +
      (src105[86] << 105) +
      (src105[87] << 105) +
      (src105[88] << 105) +
      (src105[89] << 105) +
      (src105[90] << 105) +
      (src105[91] << 105) +
      (src105[92] << 105) +
      (src105[93] << 105) +
      (src105[94] << 105) +
      (src105[95] << 105) +
      (src105[96] << 105) +
      (src105[97] << 105) +
      (src105[98] << 105) +
      (src105[99] << 105) +
      (src105[100] << 105) +
      (src105[101] << 105) +
      (src105[102] << 105) +
      (src105[103] << 105) +
      (src105[104] << 105) +
      (src105[105] << 105) +
      (src105[106] << 105) +
      (src105[107] << 105) +
      (src105[108] << 105) +
      (src105[109] << 105) +
      (src105[110] << 105) +
      (src105[111] << 105) +
      (src105[112] << 105) +
      (src105[113] << 105) +
      (src105[114] << 105) +
      (src105[115] << 105) +
      (src105[116] << 105) +
      (src105[117] << 105) +
      (src105[118] << 105) +
      (src105[119] << 105) +
      (src105[120] << 105) +
      (src105[121] << 105) +
      (src105[122] << 105) +
      (src105[123] << 105) +
      (src105[124] << 105) +
      (src105[125] << 105) +
      (src105[126] << 105) +
      (src105[127] << 105) +
      (src106[0] << 106) +
      (src106[1] << 106) +
      (src106[2] << 106) +
      (src106[3] << 106) +
      (src106[4] << 106) +
      (src106[5] << 106) +
      (src106[6] << 106) +
      (src106[7] << 106) +
      (src106[8] << 106) +
      (src106[9] << 106) +
      (src106[10] << 106) +
      (src106[11] << 106) +
      (src106[12] << 106) +
      (src106[13] << 106) +
      (src106[14] << 106) +
      (src106[15] << 106) +
      (src106[16] << 106) +
      (src106[17] << 106) +
      (src106[18] << 106) +
      (src106[19] << 106) +
      (src106[20] << 106) +
      (src106[21] << 106) +
      (src106[22] << 106) +
      (src106[23] << 106) +
      (src106[24] << 106) +
      (src106[25] << 106) +
      (src106[26] << 106) +
      (src106[27] << 106) +
      (src106[28] << 106) +
      (src106[29] << 106) +
      (src106[30] << 106) +
      (src106[31] << 106) +
      (src106[32] << 106) +
      (src106[33] << 106) +
      (src106[34] << 106) +
      (src106[35] << 106) +
      (src106[36] << 106) +
      (src106[37] << 106) +
      (src106[38] << 106) +
      (src106[39] << 106) +
      (src106[40] << 106) +
      (src106[41] << 106) +
      (src106[42] << 106) +
      (src106[43] << 106) +
      (src106[44] << 106) +
      (src106[45] << 106) +
      (src106[46] << 106) +
      (src106[47] << 106) +
      (src106[48] << 106) +
      (src106[49] << 106) +
      (src106[50] << 106) +
      (src106[51] << 106) +
      (src106[52] << 106) +
      (src106[53] << 106) +
      (src106[54] << 106) +
      (src106[55] << 106) +
      (src106[56] << 106) +
      (src106[57] << 106) +
      (src106[58] << 106) +
      (src106[59] << 106) +
      (src106[60] << 106) +
      (src106[61] << 106) +
      (src106[62] << 106) +
      (src106[63] << 106) +
      (src106[64] << 106) +
      (src106[65] << 106) +
      (src106[66] << 106) +
      (src106[67] << 106) +
      (src106[68] << 106) +
      (src106[69] << 106) +
      (src106[70] << 106) +
      (src106[71] << 106) +
      (src106[72] << 106) +
      (src106[73] << 106) +
      (src106[74] << 106) +
      (src106[75] << 106) +
      (src106[76] << 106) +
      (src106[77] << 106) +
      (src106[78] << 106) +
      (src106[79] << 106) +
      (src106[80] << 106) +
      (src106[81] << 106) +
      (src106[82] << 106) +
      (src106[83] << 106) +
      (src106[84] << 106) +
      (src106[85] << 106) +
      (src106[86] << 106) +
      (src106[87] << 106) +
      (src106[88] << 106) +
      (src106[89] << 106) +
      (src106[90] << 106) +
      (src106[91] << 106) +
      (src106[92] << 106) +
      (src106[93] << 106) +
      (src106[94] << 106) +
      (src106[95] << 106) +
      (src106[96] << 106) +
      (src106[97] << 106) +
      (src106[98] << 106) +
      (src106[99] << 106) +
      (src106[100] << 106) +
      (src106[101] << 106) +
      (src106[102] << 106) +
      (src106[103] << 106) +
      (src106[104] << 106) +
      (src106[105] << 106) +
      (src106[106] << 106) +
      (src106[107] << 106) +
      (src106[108] << 106) +
      (src106[109] << 106) +
      (src106[110] << 106) +
      (src106[111] << 106) +
      (src106[112] << 106) +
      (src106[113] << 106) +
      (src106[114] << 106) +
      (src106[115] << 106) +
      (src106[116] << 106) +
      (src106[117] << 106) +
      (src106[118] << 106) +
      (src106[119] << 106) +
      (src106[120] << 106) +
      (src106[121] << 106) +
      (src106[122] << 106) +
      (src106[123] << 106) +
      (src106[124] << 106) +
      (src106[125] << 106) +
      (src106[126] << 106) +
      (src106[127] << 106) +
      (src107[0] << 107) +
      (src107[1] << 107) +
      (src107[2] << 107) +
      (src107[3] << 107) +
      (src107[4] << 107) +
      (src107[5] << 107) +
      (src107[6] << 107) +
      (src107[7] << 107) +
      (src107[8] << 107) +
      (src107[9] << 107) +
      (src107[10] << 107) +
      (src107[11] << 107) +
      (src107[12] << 107) +
      (src107[13] << 107) +
      (src107[14] << 107) +
      (src107[15] << 107) +
      (src107[16] << 107) +
      (src107[17] << 107) +
      (src107[18] << 107) +
      (src107[19] << 107) +
      (src107[20] << 107) +
      (src107[21] << 107) +
      (src107[22] << 107) +
      (src107[23] << 107) +
      (src107[24] << 107) +
      (src107[25] << 107) +
      (src107[26] << 107) +
      (src107[27] << 107) +
      (src107[28] << 107) +
      (src107[29] << 107) +
      (src107[30] << 107) +
      (src107[31] << 107) +
      (src107[32] << 107) +
      (src107[33] << 107) +
      (src107[34] << 107) +
      (src107[35] << 107) +
      (src107[36] << 107) +
      (src107[37] << 107) +
      (src107[38] << 107) +
      (src107[39] << 107) +
      (src107[40] << 107) +
      (src107[41] << 107) +
      (src107[42] << 107) +
      (src107[43] << 107) +
      (src107[44] << 107) +
      (src107[45] << 107) +
      (src107[46] << 107) +
      (src107[47] << 107) +
      (src107[48] << 107) +
      (src107[49] << 107) +
      (src107[50] << 107) +
      (src107[51] << 107) +
      (src107[52] << 107) +
      (src107[53] << 107) +
      (src107[54] << 107) +
      (src107[55] << 107) +
      (src107[56] << 107) +
      (src107[57] << 107) +
      (src107[58] << 107) +
      (src107[59] << 107) +
      (src107[60] << 107) +
      (src107[61] << 107) +
      (src107[62] << 107) +
      (src107[63] << 107) +
      (src107[64] << 107) +
      (src107[65] << 107) +
      (src107[66] << 107) +
      (src107[67] << 107) +
      (src107[68] << 107) +
      (src107[69] << 107) +
      (src107[70] << 107) +
      (src107[71] << 107) +
      (src107[72] << 107) +
      (src107[73] << 107) +
      (src107[74] << 107) +
      (src107[75] << 107) +
      (src107[76] << 107) +
      (src107[77] << 107) +
      (src107[78] << 107) +
      (src107[79] << 107) +
      (src107[80] << 107) +
      (src107[81] << 107) +
      (src107[82] << 107) +
      (src107[83] << 107) +
      (src107[84] << 107) +
      (src107[85] << 107) +
      (src107[86] << 107) +
      (src107[87] << 107) +
      (src107[88] << 107) +
      (src107[89] << 107) +
      (src107[90] << 107) +
      (src107[91] << 107) +
      (src107[92] << 107) +
      (src107[93] << 107) +
      (src107[94] << 107) +
      (src107[95] << 107) +
      (src107[96] << 107) +
      (src107[97] << 107) +
      (src107[98] << 107) +
      (src107[99] << 107) +
      (src107[100] << 107) +
      (src107[101] << 107) +
      (src107[102] << 107) +
      (src107[103] << 107) +
      (src107[104] << 107) +
      (src107[105] << 107) +
      (src107[106] << 107) +
      (src107[107] << 107) +
      (src107[108] << 107) +
      (src107[109] << 107) +
      (src107[110] << 107) +
      (src107[111] << 107) +
      (src107[112] << 107) +
      (src107[113] << 107) +
      (src107[114] << 107) +
      (src107[115] << 107) +
      (src107[116] << 107) +
      (src107[117] << 107) +
      (src107[118] << 107) +
      (src107[119] << 107) +
      (src107[120] << 107) +
      (src107[121] << 107) +
      (src107[122] << 107) +
      (src107[123] << 107) +
      (src107[124] << 107) +
      (src107[125] << 107) +
      (src107[126] << 107) +
      (src107[127] << 107) +
      (src108[0] << 108) +
      (src108[1] << 108) +
      (src108[2] << 108) +
      (src108[3] << 108) +
      (src108[4] << 108) +
      (src108[5] << 108) +
      (src108[6] << 108) +
      (src108[7] << 108) +
      (src108[8] << 108) +
      (src108[9] << 108) +
      (src108[10] << 108) +
      (src108[11] << 108) +
      (src108[12] << 108) +
      (src108[13] << 108) +
      (src108[14] << 108) +
      (src108[15] << 108) +
      (src108[16] << 108) +
      (src108[17] << 108) +
      (src108[18] << 108) +
      (src108[19] << 108) +
      (src108[20] << 108) +
      (src108[21] << 108) +
      (src108[22] << 108) +
      (src108[23] << 108) +
      (src108[24] << 108) +
      (src108[25] << 108) +
      (src108[26] << 108) +
      (src108[27] << 108) +
      (src108[28] << 108) +
      (src108[29] << 108) +
      (src108[30] << 108) +
      (src108[31] << 108) +
      (src108[32] << 108) +
      (src108[33] << 108) +
      (src108[34] << 108) +
      (src108[35] << 108) +
      (src108[36] << 108) +
      (src108[37] << 108) +
      (src108[38] << 108) +
      (src108[39] << 108) +
      (src108[40] << 108) +
      (src108[41] << 108) +
      (src108[42] << 108) +
      (src108[43] << 108) +
      (src108[44] << 108) +
      (src108[45] << 108) +
      (src108[46] << 108) +
      (src108[47] << 108) +
      (src108[48] << 108) +
      (src108[49] << 108) +
      (src108[50] << 108) +
      (src108[51] << 108) +
      (src108[52] << 108) +
      (src108[53] << 108) +
      (src108[54] << 108) +
      (src108[55] << 108) +
      (src108[56] << 108) +
      (src108[57] << 108) +
      (src108[58] << 108) +
      (src108[59] << 108) +
      (src108[60] << 108) +
      (src108[61] << 108) +
      (src108[62] << 108) +
      (src108[63] << 108) +
      (src108[64] << 108) +
      (src108[65] << 108) +
      (src108[66] << 108) +
      (src108[67] << 108) +
      (src108[68] << 108) +
      (src108[69] << 108) +
      (src108[70] << 108) +
      (src108[71] << 108) +
      (src108[72] << 108) +
      (src108[73] << 108) +
      (src108[74] << 108) +
      (src108[75] << 108) +
      (src108[76] << 108) +
      (src108[77] << 108) +
      (src108[78] << 108) +
      (src108[79] << 108) +
      (src108[80] << 108) +
      (src108[81] << 108) +
      (src108[82] << 108) +
      (src108[83] << 108) +
      (src108[84] << 108) +
      (src108[85] << 108) +
      (src108[86] << 108) +
      (src108[87] << 108) +
      (src108[88] << 108) +
      (src108[89] << 108) +
      (src108[90] << 108) +
      (src108[91] << 108) +
      (src108[92] << 108) +
      (src108[93] << 108) +
      (src108[94] << 108) +
      (src108[95] << 108) +
      (src108[96] << 108) +
      (src108[97] << 108) +
      (src108[98] << 108) +
      (src108[99] << 108) +
      (src108[100] << 108) +
      (src108[101] << 108) +
      (src108[102] << 108) +
      (src108[103] << 108) +
      (src108[104] << 108) +
      (src108[105] << 108) +
      (src108[106] << 108) +
      (src108[107] << 108) +
      (src108[108] << 108) +
      (src108[109] << 108) +
      (src108[110] << 108) +
      (src108[111] << 108) +
      (src108[112] << 108) +
      (src108[113] << 108) +
      (src108[114] << 108) +
      (src108[115] << 108) +
      (src108[116] << 108) +
      (src108[117] << 108) +
      (src108[118] << 108) +
      (src108[119] << 108) +
      (src108[120] << 108) +
      (src108[121] << 108) +
      (src108[122] << 108) +
      (src108[123] << 108) +
      (src108[124] << 108) +
      (src108[125] << 108) +
      (src108[126] << 108) +
      (src108[127] << 108) +
      (src109[0] << 109) +
      (src109[1] << 109) +
      (src109[2] << 109) +
      (src109[3] << 109) +
      (src109[4] << 109) +
      (src109[5] << 109) +
      (src109[6] << 109) +
      (src109[7] << 109) +
      (src109[8] << 109) +
      (src109[9] << 109) +
      (src109[10] << 109) +
      (src109[11] << 109) +
      (src109[12] << 109) +
      (src109[13] << 109) +
      (src109[14] << 109) +
      (src109[15] << 109) +
      (src109[16] << 109) +
      (src109[17] << 109) +
      (src109[18] << 109) +
      (src109[19] << 109) +
      (src109[20] << 109) +
      (src109[21] << 109) +
      (src109[22] << 109) +
      (src109[23] << 109) +
      (src109[24] << 109) +
      (src109[25] << 109) +
      (src109[26] << 109) +
      (src109[27] << 109) +
      (src109[28] << 109) +
      (src109[29] << 109) +
      (src109[30] << 109) +
      (src109[31] << 109) +
      (src109[32] << 109) +
      (src109[33] << 109) +
      (src109[34] << 109) +
      (src109[35] << 109) +
      (src109[36] << 109) +
      (src109[37] << 109) +
      (src109[38] << 109) +
      (src109[39] << 109) +
      (src109[40] << 109) +
      (src109[41] << 109) +
      (src109[42] << 109) +
      (src109[43] << 109) +
      (src109[44] << 109) +
      (src109[45] << 109) +
      (src109[46] << 109) +
      (src109[47] << 109) +
      (src109[48] << 109) +
      (src109[49] << 109) +
      (src109[50] << 109) +
      (src109[51] << 109) +
      (src109[52] << 109) +
      (src109[53] << 109) +
      (src109[54] << 109) +
      (src109[55] << 109) +
      (src109[56] << 109) +
      (src109[57] << 109) +
      (src109[58] << 109) +
      (src109[59] << 109) +
      (src109[60] << 109) +
      (src109[61] << 109) +
      (src109[62] << 109) +
      (src109[63] << 109) +
      (src109[64] << 109) +
      (src109[65] << 109) +
      (src109[66] << 109) +
      (src109[67] << 109) +
      (src109[68] << 109) +
      (src109[69] << 109) +
      (src109[70] << 109) +
      (src109[71] << 109) +
      (src109[72] << 109) +
      (src109[73] << 109) +
      (src109[74] << 109) +
      (src109[75] << 109) +
      (src109[76] << 109) +
      (src109[77] << 109) +
      (src109[78] << 109) +
      (src109[79] << 109) +
      (src109[80] << 109) +
      (src109[81] << 109) +
      (src109[82] << 109) +
      (src109[83] << 109) +
      (src109[84] << 109) +
      (src109[85] << 109) +
      (src109[86] << 109) +
      (src109[87] << 109) +
      (src109[88] << 109) +
      (src109[89] << 109) +
      (src109[90] << 109) +
      (src109[91] << 109) +
      (src109[92] << 109) +
      (src109[93] << 109) +
      (src109[94] << 109) +
      (src109[95] << 109) +
      (src109[96] << 109) +
      (src109[97] << 109) +
      (src109[98] << 109) +
      (src109[99] << 109) +
      (src109[100] << 109) +
      (src109[101] << 109) +
      (src109[102] << 109) +
      (src109[103] << 109) +
      (src109[104] << 109) +
      (src109[105] << 109) +
      (src109[106] << 109) +
      (src109[107] << 109) +
      (src109[108] << 109) +
      (src109[109] << 109) +
      (src109[110] << 109) +
      (src109[111] << 109) +
      (src109[112] << 109) +
      (src109[113] << 109) +
      (src109[114] << 109) +
      (src109[115] << 109) +
      (src109[116] << 109) +
      (src109[117] << 109) +
      (src109[118] << 109) +
      (src109[119] << 109) +
      (src109[120] << 109) +
      (src109[121] << 109) +
      (src109[122] << 109) +
      (src109[123] << 109) +
      (src109[124] << 109) +
      (src109[125] << 109) +
      (src109[126] << 109) +
      (src109[127] << 109) +
      (src110[0] << 110) +
      (src110[1] << 110) +
      (src110[2] << 110) +
      (src110[3] << 110) +
      (src110[4] << 110) +
      (src110[5] << 110) +
      (src110[6] << 110) +
      (src110[7] << 110) +
      (src110[8] << 110) +
      (src110[9] << 110) +
      (src110[10] << 110) +
      (src110[11] << 110) +
      (src110[12] << 110) +
      (src110[13] << 110) +
      (src110[14] << 110) +
      (src110[15] << 110) +
      (src110[16] << 110) +
      (src110[17] << 110) +
      (src110[18] << 110) +
      (src110[19] << 110) +
      (src110[20] << 110) +
      (src110[21] << 110) +
      (src110[22] << 110) +
      (src110[23] << 110) +
      (src110[24] << 110) +
      (src110[25] << 110) +
      (src110[26] << 110) +
      (src110[27] << 110) +
      (src110[28] << 110) +
      (src110[29] << 110) +
      (src110[30] << 110) +
      (src110[31] << 110) +
      (src110[32] << 110) +
      (src110[33] << 110) +
      (src110[34] << 110) +
      (src110[35] << 110) +
      (src110[36] << 110) +
      (src110[37] << 110) +
      (src110[38] << 110) +
      (src110[39] << 110) +
      (src110[40] << 110) +
      (src110[41] << 110) +
      (src110[42] << 110) +
      (src110[43] << 110) +
      (src110[44] << 110) +
      (src110[45] << 110) +
      (src110[46] << 110) +
      (src110[47] << 110) +
      (src110[48] << 110) +
      (src110[49] << 110) +
      (src110[50] << 110) +
      (src110[51] << 110) +
      (src110[52] << 110) +
      (src110[53] << 110) +
      (src110[54] << 110) +
      (src110[55] << 110) +
      (src110[56] << 110) +
      (src110[57] << 110) +
      (src110[58] << 110) +
      (src110[59] << 110) +
      (src110[60] << 110) +
      (src110[61] << 110) +
      (src110[62] << 110) +
      (src110[63] << 110) +
      (src110[64] << 110) +
      (src110[65] << 110) +
      (src110[66] << 110) +
      (src110[67] << 110) +
      (src110[68] << 110) +
      (src110[69] << 110) +
      (src110[70] << 110) +
      (src110[71] << 110) +
      (src110[72] << 110) +
      (src110[73] << 110) +
      (src110[74] << 110) +
      (src110[75] << 110) +
      (src110[76] << 110) +
      (src110[77] << 110) +
      (src110[78] << 110) +
      (src110[79] << 110) +
      (src110[80] << 110) +
      (src110[81] << 110) +
      (src110[82] << 110) +
      (src110[83] << 110) +
      (src110[84] << 110) +
      (src110[85] << 110) +
      (src110[86] << 110) +
      (src110[87] << 110) +
      (src110[88] << 110) +
      (src110[89] << 110) +
      (src110[90] << 110) +
      (src110[91] << 110) +
      (src110[92] << 110) +
      (src110[93] << 110) +
      (src110[94] << 110) +
      (src110[95] << 110) +
      (src110[96] << 110) +
      (src110[97] << 110) +
      (src110[98] << 110) +
      (src110[99] << 110) +
      (src110[100] << 110) +
      (src110[101] << 110) +
      (src110[102] << 110) +
      (src110[103] << 110) +
      (src110[104] << 110) +
      (src110[105] << 110) +
      (src110[106] << 110) +
      (src110[107] << 110) +
      (src110[108] << 110) +
      (src110[109] << 110) +
      (src110[110] << 110) +
      (src110[111] << 110) +
      (src110[112] << 110) +
      (src110[113] << 110) +
      (src110[114] << 110) +
      (src110[115] << 110) +
      (src110[116] << 110) +
      (src110[117] << 110) +
      (src110[118] << 110) +
      (src110[119] << 110) +
      (src110[120] << 110) +
      (src110[121] << 110) +
      (src110[122] << 110) +
      (src110[123] << 110) +
      (src110[124] << 110) +
      (src110[125] << 110) +
      (src110[126] << 110) +
      (src110[127] << 110) +
      (src111[0] << 111) +
      (src111[1] << 111) +
      (src111[2] << 111) +
      (src111[3] << 111) +
      (src111[4] << 111) +
      (src111[5] << 111) +
      (src111[6] << 111) +
      (src111[7] << 111) +
      (src111[8] << 111) +
      (src111[9] << 111) +
      (src111[10] << 111) +
      (src111[11] << 111) +
      (src111[12] << 111) +
      (src111[13] << 111) +
      (src111[14] << 111) +
      (src111[15] << 111) +
      (src111[16] << 111) +
      (src111[17] << 111) +
      (src111[18] << 111) +
      (src111[19] << 111) +
      (src111[20] << 111) +
      (src111[21] << 111) +
      (src111[22] << 111) +
      (src111[23] << 111) +
      (src111[24] << 111) +
      (src111[25] << 111) +
      (src111[26] << 111) +
      (src111[27] << 111) +
      (src111[28] << 111) +
      (src111[29] << 111) +
      (src111[30] << 111) +
      (src111[31] << 111) +
      (src111[32] << 111) +
      (src111[33] << 111) +
      (src111[34] << 111) +
      (src111[35] << 111) +
      (src111[36] << 111) +
      (src111[37] << 111) +
      (src111[38] << 111) +
      (src111[39] << 111) +
      (src111[40] << 111) +
      (src111[41] << 111) +
      (src111[42] << 111) +
      (src111[43] << 111) +
      (src111[44] << 111) +
      (src111[45] << 111) +
      (src111[46] << 111) +
      (src111[47] << 111) +
      (src111[48] << 111) +
      (src111[49] << 111) +
      (src111[50] << 111) +
      (src111[51] << 111) +
      (src111[52] << 111) +
      (src111[53] << 111) +
      (src111[54] << 111) +
      (src111[55] << 111) +
      (src111[56] << 111) +
      (src111[57] << 111) +
      (src111[58] << 111) +
      (src111[59] << 111) +
      (src111[60] << 111) +
      (src111[61] << 111) +
      (src111[62] << 111) +
      (src111[63] << 111) +
      (src111[64] << 111) +
      (src111[65] << 111) +
      (src111[66] << 111) +
      (src111[67] << 111) +
      (src111[68] << 111) +
      (src111[69] << 111) +
      (src111[70] << 111) +
      (src111[71] << 111) +
      (src111[72] << 111) +
      (src111[73] << 111) +
      (src111[74] << 111) +
      (src111[75] << 111) +
      (src111[76] << 111) +
      (src111[77] << 111) +
      (src111[78] << 111) +
      (src111[79] << 111) +
      (src111[80] << 111) +
      (src111[81] << 111) +
      (src111[82] << 111) +
      (src111[83] << 111) +
      (src111[84] << 111) +
      (src111[85] << 111) +
      (src111[86] << 111) +
      (src111[87] << 111) +
      (src111[88] << 111) +
      (src111[89] << 111) +
      (src111[90] << 111) +
      (src111[91] << 111) +
      (src111[92] << 111) +
      (src111[93] << 111) +
      (src111[94] << 111) +
      (src111[95] << 111) +
      (src111[96] << 111) +
      (src111[97] << 111) +
      (src111[98] << 111) +
      (src111[99] << 111) +
      (src111[100] << 111) +
      (src111[101] << 111) +
      (src111[102] << 111) +
      (src111[103] << 111) +
      (src111[104] << 111) +
      (src111[105] << 111) +
      (src111[106] << 111) +
      (src111[107] << 111) +
      (src111[108] << 111) +
      (src111[109] << 111) +
      (src111[110] << 111) +
      (src111[111] << 111) +
      (src111[112] << 111) +
      (src111[113] << 111) +
      (src111[114] << 111) +
      (src111[115] << 111) +
      (src111[116] << 111) +
      (src111[117] << 111) +
      (src111[118] << 111) +
      (src111[119] << 111) +
      (src111[120] << 111) +
      (src111[121] << 111) +
      (src111[122] << 111) +
      (src111[123] << 111) +
      (src111[124] << 111) +
      (src111[125] << 111) +
      (src111[126] << 111) +
      (src111[127] << 111) +
      (src112[0] << 112) +
      (src112[1] << 112) +
      (src112[2] << 112) +
      (src112[3] << 112) +
      (src112[4] << 112) +
      (src112[5] << 112) +
      (src112[6] << 112) +
      (src112[7] << 112) +
      (src112[8] << 112) +
      (src112[9] << 112) +
      (src112[10] << 112) +
      (src112[11] << 112) +
      (src112[12] << 112) +
      (src112[13] << 112) +
      (src112[14] << 112) +
      (src112[15] << 112) +
      (src112[16] << 112) +
      (src112[17] << 112) +
      (src112[18] << 112) +
      (src112[19] << 112) +
      (src112[20] << 112) +
      (src112[21] << 112) +
      (src112[22] << 112) +
      (src112[23] << 112) +
      (src112[24] << 112) +
      (src112[25] << 112) +
      (src112[26] << 112) +
      (src112[27] << 112) +
      (src112[28] << 112) +
      (src112[29] << 112) +
      (src112[30] << 112) +
      (src112[31] << 112) +
      (src112[32] << 112) +
      (src112[33] << 112) +
      (src112[34] << 112) +
      (src112[35] << 112) +
      (src112[36] << 112) +
      (src112[37] << 112) +
      (src112[38] << 112) +
      (src112[39] << 112) +
      (src112[40] << 112) +
      (src112[41] << 112) +
      (src112[42] << 112) +
      (src112[43] << 112) +
      (src112[44] << 112) +
      (src112[45] << 112) +
      (src112[46] << 112) +
      (src112[47] << 112) +
      (src112[48] << 112) +
      (src112[49] << 112) +
      (src112[50] << 112) +
      (src112[51] << 112) +
      (src112[52] << 112) +
      (src112[53] << 112) +
      (src112[54] << 112) +
      (src112[55] << 112) +
      (src112[56] << 112) +
      (src112[57] << 112) +
      (src112[58] << 112) +
      (src112[59] << 112) +
      (src112[60] << 112) +
      (src112[61] << 112) +
      (src112[62] << 112) +
      (src112[63] << 112) +
      (src112[64] << 112) +
      (src112[65] << 112) +
      (src112[66] << 112) +
      (src112[67] << 112) +
      (src112[68] << 112) +
      (src112[69] << 112) +
      (src112[70] << 112) +
      (src112[71] << 112) +
      (src112[72] << 112) +
      (src112[73] << 112) +
      (src112[74] << 112) +
      (src112[75] << 112) +
      (src112[76] << 112) +
      (src112[77] << 112) +
      (src112[78] << 112) +
      (src112[79] << 112) +
      (src112[80] << 112) +
      (src112[81] << 112) +
      (src112[82] << 112) +
      (src112[83] << 112) +
      (src112[84] << 112) +
      (src112[85] << 112) +
      (src112[86] << 112) +
      (src112[87] << 112) +
      (src112[88] << 112) +
      (src112[89] << 112) +
      (src112[90] << 112) +
      (src112[91] << 112) +
      (src112[92] << 112) +
      (src112[93] << 112) +
      (src112[94] << 112) +
      (src112[95] << 112) +
      (src112[96] << 112) +
      (src112[97] << 112) +
      (src112[98] << 112) +
      (src112[99] << 112) +
      (src112[100] << 112) +
      (src112[101] << 112) +
      (src112[102] << 112) +
      (src112[103] << 112) +
      (src112[104] << 112) +
      (src112[105] << 112) +
      (src112[106] << 112) +
      (src112[107] << 112) +
      (src112[108] << 112) +
      (src112[109] << 112) +
      (src112[110] << 112) +
      (src112[111] << 112) +
      (src112[112] << 112) +
      (src112[113] << 112) +
      (src112[114] << 112) +
      (src112[115] << 112) +
      (src112[116] << 112) +
      (src112[117] << 112) +
      (src112[118] << 112) +
      (src112[119] << 112) +
      (src112[120] << 112) +
      (src112[121] << 112) +
      (src112[122] << 112) +
      (src112[123] << 112) +
      (src112[124] << 112) +
      (src112[125] << 112) +
      (src112[126] << 112) +
      (src112[127] << 112) +
      (src113[0] << 113) +
      (src113[1] << 113) +
      (src113[2] << 113) +
      (src113[3] << 113) +
      (src113[4] << 113) +
      (src113[5] << 113) +
      (src113[6] << 113) +
      (src113[7] << 113) +
      (src113[8] << 113) +
      (src113[9] << 113) +
      (src113[10] << 113) +
      (src113[11] << 113) +
      (src113[12] << 113) +
      (src113[13] << 113) +
      (src113[14] << 113) +
      (src113[15] << 113) +
      (src113[16] << 113) +
      (src113[17] << 113) +
      (src113[18] << 113) +
      (src113[19] << 113) +
      (src113[20] << 113) +
      (src113[21] << 113) +
      (src113[22] << 113) +
      (src113[23] << 113) +
      (src113[24] << 113) +
      (src113[25] << 113) +
      (src113[26] << 113) +
      (src113[27] << 113) +
      (src113[28] << 113) +
      (src113[29] << 113) +
      (src113[30] << 113) +
      (src113[31] << 113) +
      (src113[32] << 113) +
      (src113[33] << 113) +
      (src113[34] << 113) +
      (src113[35] << 113) +
      (src113[36] << 113) +
      (src113[37] << 113) +
      (src113[38] << 113) +
      (src113[39] << 113) +
      (src113[40] << 113) +
      (src113[41] << 113) +
      (src113[42] << 113) +
      (src113[43] << 113) +
      (src113[44] << 113) +
      (src113[45] << 113) +
      (src113[46] << 113) +
      (src113[47] << 113) +
      (src113[48] << 113) +
      (src113[49] << 113) +
      (src113[50] << 113) +
      (src113[51] << 113) +
      (src113[52] << 113) +
      (src113[53] << 113) +
      (src113[54] << 113) +
      (src113[55] << 113) +
      (src113[56] << 113) +
      (src113[57] << 113) +
      (src113[58] << 113) +
      (src113[59] << 113) +
      (src113[60] << 113) +
      (src113[61] << 113) +
      (src113[62] << 113) +
      (src113[63] << 113) +
      (src113[64] << 113) +
      (src113[65] << 113) +
      (src113[66] << 113) +
      (src113[67] << 113) +
      (src113[68] << 113) +
      (src113[69] << 113) +
      (src113[70] << 113) +
      (src113[71] << 113) +
      (src113[72] << 113) +
      (src113[73] << 113) +
      (src113[74] << 113) +
      (src113[75] << 113) +
      (src113[76] << 113) +
      (src113[77] << 113) +
      (src113[78] << 113) +
      (src113[79] << 113) +
      (src113[80] << 113) +
      (src113[81] << 113) +
      (src113[82] << 113) +
      (src113[83] << 113) +
      (src113[84] << 113) +
      (src113[85] << 113) +
      (src113[86] << 113) +
      (src113[87] << 113) +
      (src113[88] << 113) +
      (src113[89] << 113) +
      (src113[90] << 113) +
      (src113[91] << 113) +
      (src113[92] << 113) +
      (src113[93] << 113) +
      (src113[94] << 113) +
      (src113[95] << 113) +
      (src113[96] << 113) +
      (src113[97] << 113) +
      (src113[98] << 113) +
      (src113[99] << 113) +
      (src113[100] << 113) +
      (src113[101] << 113) +
      (src113[102] << 113) +
      (src113[103] << 113) +
      (src113[104] << 113) +
      (src113[105] << 113) +
      (src113[106] << 113) +
      (src113[107] << 113) +
      (src113[108] << 113) +
      (src113[109] << 113) +
      (src113[110] << 113) +
      (src113[111] << 113) +
      (src113[112] << 113) +
      (src113[113] << 113) +
      (src113[114] << 113) +
      (src113[115] << 113) +
      (src113[116] << 113) +
      (src113[117] << 113) +
      (src113[118] << 113) +
      (src113[119] << 113) +
      (src113[120] << 113) +
      (src113[121] << 113) +
      (src113[122] << 113) +
      (src113[123] << 113) +
      (src113[124] << 113) +
      (src113[125] << 113) +
      (src113[126] << 113) +
      (src113[127] << 113) +
      (src114[0] << 114) +
      (src114[1] << 114) +
      (src114[2] << 114) +
      (src114[3] << 114) +
      (src114[4] << 114) +
      (src114[5] << 114) +
      (src114[6] << 114) +
      (src114[7] << 114) +
      (src114[8] << 114) +
      (src114[9] << 114) +
      (src114[10] << 114) +
      (src114[11] << 114) +
      (src114[12] << 114) +
      (src114[13] << 114) +
      (src114[14] << 114) +
      (src114[15] << 114) +
      (src114[16] << 114) +
      (src114[17] << 114) +
      (src114[18] << 114) +
      (src114[19] << 114) +
      (src114[20] << 114) +
      (src114[21] << 114) +
      (src114[22] << 114) +
      (src114[23] << 114) +
      (src114[24] << 114) +
      (src114[25] << 114) +
      (src114[26] << 114) +
      (src114[27] << 114) +
      (src114[28] << 114) +
      (src114[29] << 114) +
      (src114[30] << 114) +
      (src114[31] << 114) +
      (src114[32] << 114) +
      (src114[33] << 114) +
      (src114[34] << 114) +
      (src114[35] << 114) +
      (src114[36] << 114) +
      (src114[37] << 114) +
      (src114[38] << 114) +
      (src114[39] << 114) +
      (src114[40] << 114) +
      (src114[41] << 114) +
      (src114[42] << 114) +
      (src114[43] << 114) +
      (src114[44] << 114) +
      (src114[45] << 114) +
      (src114[46] << 114) +
      (src114[47] << 114) +
      (src114[48] << 114) +
      (src114[49] << 114) +
      (src114[50] << 114) +
      (src114[51] << 114) +
      (src114[52] << 114) +
      (src114[53] << 114) +
      (src114[54] << 114) +
      (src114[55] << 114) +
      (src114[56] << 114) +
      (src114[57] << 114) +
      (src114[58] << 114) +
      (src114[59] << 114) +
      (src114[60] << 114) +
      (src114[61] << 114) +
      (src114[62] << 114) +
      (src114[63] << 114) +
      (src114[64] << 114) +
      (src114[65] << 114) +
      (src114[66] << 114) +
      (src114[67] << 114) +
      (src114[68] << 114) +
      (src114[69] << 114) +
      (src114[70] << 114) +
      (src114[71] << 114) +
      (src114[72] << 114) +
      (src114[73] << 114) +
      (src114[74] << 114) +
      (src114[75] << 114) +
      (src114[76] << 114) +
      (src114[77] << 114) +
      (src114[78] << 114) +
      (src114[79] << 114) +
      (src114[80] << 114) +
      (src114[81] << 114) +
      (src114[82] << 114) +
      (src114[83] << 114) +
      (src114[84] << 114) +
      (src114[85] << 114) +
      (src114[86] << 114) +
      (src114[87] << 114) +
      (src114[88] << 114) +
      (src114[89] << 114) +
      (src114[90] << 114) +
      (src114[91] << 114) +
      (src114[92] << 114) +
      (src114[93] << 114) +
      (src114[94] << 114) +
      (src114[95] << 114) +
      (src114[96] << 114) +
      (src114[97] << 114) +
      (src114[98] << 114) +
      (src114[99] << 114) +
      (src114[100] << 114) +
      (src114[101] << 114) +
      (src114[102] << 114) +
      (src114[103] << 114) +
      (src114[104] << 114) +
      (src114[105] << 114) +
      (src114[106] << 114) +
      (src114[107] << 114) +
      (src114[108] << 114) +
      (src114[109] << 114) +
      (src114[110] << 114) +
      (src114[111] << 114) +
      (src114[112] << 114) +
      (src114[113] << 114) +
      (src114[114] << 114) +
      (src114[115] << 114) +
      (src114[116] << 114) +
      (src114[117] << 114) +
      (src114[118] << 114) +
      (src114[119] << 114) +
      (src114[120] << 114) +
      (src114[121] << 114) +
      (src114[122] << 114) +
      (src114[123] << 114) +
      (src114[124] << 114) +
      (src114[125] << 114) +
      (src114[126] << 114) +
      (src114[127] << 114) +
      (src115[0] << 115) +
      (src115[1] << 115) +
      (src115[2] << 115) +
      (src115[3] << 115) +
      (src115[4] << 115) +
      (src115[5] << 115) +
      (src115[6] << 115) +
      (src115[7] << 115) +
      (src115[8] << 115) +
      (src115[9] << 115) +
      (src115[10] << 115) +
      (src115[11] << 115) +
      (src115[12] << 115) +
      (src115[13] << 115) +
      (src115[14] << 115) +
      (src115[15] << 115) +
      (src115[16] << 115) +
      (src115[17] << 115) +
      (src115[18] << 115) +
      (src115[19] << 115) +
      (src115[20] << 115) +
      (src115[21] << 115) +
      (src115[22] << 115) +
      (src115[23] << 115) +
      (src115[24] << 115) +
      (src115[25] << 115) +
      (src115[26] << 115) +
      (src115[27] << 115) +
      (src115[28] << 115) +
      (src115[29] << 115) +
      (src115[30] << 115) +
      (src115[31] << 115) +
      (src115[32] << 115) +
      (src115[33] << 115) +
      (src115[34] << 115) +
      (src115[35] << 115) +
      (src115[36] << 115) +
      (src115[37] << 115) +
      (src115[38] << 115) +
      (src115[39] << 115) +
      (src115[40] << 115) +
      (src115[41] << 115) +
      (src115[42] << 115) +
      (src115[43] << 115) +
      (src115[44] << 115) +
      (src115[45] << 115) +
      (src115[46] << 115) +
      (src115[47] << 115) +
      (src115[48] << 115) +
      (src115[49] << 115) +
      (src115[50] << 115) +
      (src115[51] << 115) +
      (src115[52] << 115) +
      (src115[53] << 115) +
      (src115[54] << 115) +
      (src115[55] << 115) +
      (src115[56] << 115) +
      (src115[57] << 115) +
      (src115[58] << 115) +
      (src115[59] << 115) +
      (src115[60] << 115) +
      (src115[61] << 115) +
      (src115[62] << 115) +
      (src115[63] << 115) +
      (src115[64] << 115) +
      (src115[65] << 115) +
      (src115[66] << 115) +
      (src115[67] << 115) +
      (src115[68] << 115) +
      (src115[69] << 115) +
      (src115[70] << 115) +
      (src115[71] << 115) +
      (src115[72] << 115) +
      (src115[73] << 115) +
      (src115[74] << 115) +
      (src115[75] << 115) +
      (src115[76] << 115) +
      (src115[77] << 115) +
      (src115[78] << 115) +
      (src115[79] << 115) +
      (src115[80] << 115) +
      (src115[81] << 115) +
      (src115[82] << 115) +
      (src115[83] << 115) +
      (src115[84] << 115) +
      (src115[85] << 115) +
      (src115[86] << 115) +
      (src115[87] << 115) +
      (src115[88] << 115) +
      (src115[89] << 115) +
      (src115[90] << 115) +
      (src115[91] << 115) +
      (src115[92] << 115) +
      (src115[93] << 115) +
      (src115[94] << 115) +
      (src115[95] << 115) +
      (src115[96] << 115) +
      (src115[97] << 115) +
      (src115[98] << 115) +
      (src115[99] << 115) +
      (src115[100] << 115) +
      (src115[101] << 115) +
      (src115[102] << 115) +
      (src115[103] << 115) +
      (src115[104] << 115) +
      (src115[105] << 115) +
      (src115[106] << 115) +
      (src115[107] << 115) +
      (src115[108] << 115) +
      (src115[109] << 115) +
      (src115[110] << 115) +
      (src115[111] << 115) +
      (src115[112] << 115) +
      (src115[113] << 115) +
      (src115[114] << 115) +
      (src115[115] << 115) +
      (src115[116] << 115) +
      (src115[117] << 115) +
      (src115[118] << 115) +
      (src115[119] << 115) +
      (src115[120] << 115) +
      (src115[121] << 115) +
      (src115[122] << 115) +
      (src115[123] << 115) +
      (src115[124] << 115) +
      (src115[125] << 115) +
      (src115[126] << 115) +
      (src115[127] << 115) +
      (src116[0] << 116) +
      (src116[1] << 116) +
      (src116[2] << 116) +
      (src116[3] << 116) +
      (src116[4] << 116) +
      (src116[5] << 116) +
      (src116[6] << 116) +
      (src116[7] << 116) +
      (src116[8] << 116) +
      (src116[9] << 116) +
      (src116[10] << 116) +
      (src116[11] << 116) +
      (src116[12] << 116) +
      (src116[13] << 116) +
      (src116[14] << 116) +
      (src116[15] << 116) +
      (src116[16] << 116) +
      (src116[17] << 116) +
      (src116[18] << 116) +
      (src116[19] << 116) +
      (src116[20] << 116) +
      (src116[21] << 116) +
      (src116[22] << 116) +
      (src116[23] << 116) +
      (src116[24] << 116) +
      (src116[25] << 116) +
      (src116[26] << 116) +
      (src116[27] << 116) +
      (src116[28] << 116) +
      (src116[29] << 116) +
      (src116[30] << 116) +
      (src116[31] << 116) +
      (src116[32] << 116) +
      (src116[33] << 116) +
      (src116[34] << 116) +
      (src116[35] << 116) +
      (src116[36] << 116) +
      (src116[37] << 116) +
      (src116[38] << 116) +
      (src116[39] << 116) +
      (src116[40] << 116) +
      (src116[41] << 116) +
      (src116[42] << 116) +
      (src116[43] << 116) +
      (src116[44] << 116) +
      (src116[45] << 116) +
      (src116[46] << 116) +
      (src116[47] << 116) +
      (src116[48] << 116) +
      (src116[49] << 116) +
      (src116[50] << 116) +
      (src116[51] << 116) +
      (src116[52] << 116) +
      (src116[53] << 116) +
      (src116[54] << 116) +
      (src116[55] << 116) +
      (src116[56] << 116) +
      (src116[57] << 116) +
      (src116[58] << 116) +
      (src116[59] << 116) +
      (src116[60] << 116) +
      (src116[61] << 116) +
      (src116[62] << 116) +
      (src116[63] << 116) +
      (src116[64] << 116) +
      (src116[65] << 116) +
      (src116[66] << 116) +
      (src116[67] << 116) +
      (src116[68] << 116) +
      (src116[69] << 116) +
      (src116[70] << 116) +
      (src116[71] << 116) +
      (src116[72] << 116) +
      (src116[73] << 116) +
      (src116[74] << 116) +
      (src116[75] << 116) +
      (src116[76] << 116) +
      (src116[77] << 116) +
      (src116[78] << 116) +
      (src116[79] << 116) +
      (src116[80] << 116) +
      (src116[81] << 116) +
      (src116[82] << 116) +
      (src116[83] << 116) +
      (src116[84] << 116) +
      (src116[85] << 116) +
      (src116[86] << 116) +
      (src116[87] << 116) +
      (src116[88] << 116) +
      (src116[89] << 116) +
      (src116[90] << 116) +
      (src116[91] << 116) +
      (src116[92] << 116) +
      (src116[93] << 116) +
      (src116[94] << 116) +
      (src116[95] << 116) +
      (src116[96] << 116) +
      (src116[97] << 116) +
      (src116[98] << 116) +
      (src116[99] << 116) +
      (src116[100] << 116) +
      (src116[101] << 116) +
      (src116[102] << 116) +
      (src116[103] << 116) +
      (src116[104] << 116) +
      (src116[105] << 116) +
      (src116[106] << 116) +
      (src116[107] << 116) +
      (src116[108] << 116) +
      (src116[109] << 116) +
      (src116[110] << 116) +
      (src116[111] << 116) +
      (src116[112] << 116) +
      (src116[113] << 116) +
      (src116[114] << 116) +
      (src116[115] << 116) +
      (src116[116] << 116) +
      (src116[117] << 116) +
      (src116[118] << 116) +
      (src116[119] << 116) +
      (src116[120] << 116) +
      (src116[121] << 116) +
      (src116[122] << 116) +
      (src116[123] << 116) +
      (src116[124] << 116) +
      (src116[125] << 116) +
      (src116[126] << 116) +
      (src116[127] << 116) +
      (src117[0] << 117) +
      (src117[1] << 117) +
      (src117[2] << 117) +
      (src117[3] << 117) +
      (src117[4] << 117) +
      (src117[5] << 117) +
      (src117[6] << 117) +
      (src117[7] << 117) +
      (src117[8] << 117) +
      (src117[9] << 117) +
      (src117[10] << 117) +
      (src117[11] << 117) +
      (src117[12] << 117) +
      (src117[13] << 117) +
      (src117[14] << 117) +
      (src117[15] << 117) +
      (src117[16] << 117) +
      (src117[17] << 117) +
      (src117[18] << 117) +
      (src117[19] << 117) +
      (src117[20] << 117) +
      (src117[21] << 117) +
      (src117[22] << 117) +
      (src117[23] << 117) +
      (src117[24] << 117) +
      (src117[25] << 117) +
      (src117[26] << 117) +
      (src117[27] << 117) +
      (src117[28] << 117) +
      (src117[29] << 117) +
      (src117[30] << 117) +
      (src117[31] << 117) +
      (src117[32] << 117) +
      (src117[33] << 117) +
      (src117[34] << 117) +
      (src117[35] << 117) +
      (src117[36] << 117) +
      (src117[37] << 117) +
      (src117[38] << 117) +
      (src117[39] << 117) +
      (src117[40] << 117) +
      (src117[41] << 117) +
      (src117[42] << 117) +
      (src117[43] << 117) +
      (src117[44] << 117) +
      (src117[45] << 117) +
      (src117[46] << 117) +
      (src117[47] << 117) +
      (src117[48] << 117) +
      (src117[49] << 117) +
      (src117[50] << 117) +
      (src117[51] << 117) +
      (src117[52] << 117) +
      (src117[53] << 117) +
      (src117[54] << 117) +
      (src117[55] << 117) +
      (src117[56] << 117) +
      (src117[57] << 117) +
      (src117[58] << 117) +
      (src117[59] << 117) +
      (src117[60] << 117) +
      (src117[61] << 117) +
      (src117[62] << 117) +
      (src117[63] << 117) +
      (src117[64] << 117) +
      (src117[65] << 117) +
      (src117[66] << 117) +
      (src117[67] << 117) +
      (src117[68] << 117) +
      (src117[69] << 117) +
      (src117[70] << 117) +
      (src117[71] << 117) +
      (src117[72] << 117) +
      (src117[73] << 117) +
      (src117[74] << 117) +
      (src117[75] << 117) +
      (src117[76] << 117) +
      (src117[77] << 117) +
      (src117[78] << 117) +
      (src117[79] << 117) +
      (src117[80] << 117) +
      (src117[81] << 117) +
      (src117[82] << 117) +
      (src117[83] << 117) +
      (src117[84] << 117) +
      (src117[85] << 117) +
      (src117[86] << 117) +
      (src117[87] << 117) +
      (src117[88] << 117) +
      (src117[89] << 117) +
      (src117[90] << 117) +
      (src117[91] << 117) +
      (src117[92] << 117) +
      (src117[93] << 117) +
      (src117[94] << 117) +
      (src117[95] << 117) +
      (src117[96] << 117) +
      (src117[97] << 117) +
      (src117[98] << 117) +
      (src117[99] << 117) +
      (src117[100] << 117) +
      (src117[101] << 117) +
      (src117[102] << 117) +
      (src117[103] << 117) +
      (src117[104] << 117) +
      (src117[105] << 117) +
      (src117[106] << 117) +
      (src117[107] << 117) +
      (src117[108] << 117) +
      (src117[109] << 117) +
      (src117[110] << 117) +
      (src117[111] << 117) +
      (src117[112] << 117) +
      (src117[113] << 117) +
      (src117[114] << 117) +
      (src117[115] << 117) +
      (src117[116] << 117) +
      (src117[117] << 117) +
      (src117[118] << 117) +
      (src117[119] << 117) +
      (src117[120] << 117) +
      (src117[121] << 117) +
      (src117[122] << 117) +
      (src117[123] << 117) +
      (src117[124] << 117) +
      (src117[125] << 117) +
      (src117[126] << 117) +
      (src117[127] << 117) +
      (src118[0] << 118) +
      (src118[1] << 118) +
      (src118[2] << 118) +
      (src118[3] << 118) +
      (src118[4] << 118) +
      (src118[5] << 118) +
      (src118[6] << 118) +
      (src118[7] << 118) +
      (src118[8] << 118) +
      (src118[9] << 118) +
      (src118[10] << 118) +
      (src118[11] << 118) +
      (src118[12] << 118) +
      (src118[13] << 118) +
      (src118[14] << 118) +
      (src118[15] << 118) +
      (src118[16] << 118) +
      (src118[17] << 118) +
      (src118[18] << 118) +
      (src118[19] << 118) +
      (src118[20] << 118) +
      (src118[21] << 118) +
      (src118[22] << 118) +
      (src118[23] << 118) +
      (src118[24] << 118) +
      (src118[25] << 118) +
      (src118[26] << 118) +
      (src118[27] << 118) +
      (src118[28] << 118) +
      (src118[29] << 118) +
      (src118[30] << 118) +
      (src118[31] << 118) +
      (src118[32] << 118) +
      (src118[33] << 118) +
      (src118[34] << 118) +
      (src118[35] << 118) +
      (src118[36] << 118) +
      (src118[37] << 118) +
      (src118[38] << 118) +
      (src118[39] << 118) +
      (src118[40] << 118) +
      (src118[41] << 118) +
      (src118[42] << 118) +
      (src118[43] << 118) +
      (src118[44] << 118) +
      (src118[45] << 118) +
      (src118[46] << 118) +
      (src118[47] << 118) +
      (src118[48] << 118) +
      (src118[49] << 118) +
      (src118[50] << 118) +
      (src118[51] << 118) +
      (src118[52] << 118) +
      (src118[53] << 118) +
      (src118[54] << 118) +
      (src118[55] << 118) +
      (src118[56] << 118) +
      (src118[57] << 118) +
      (src118[58] << 118) +
      (src118[59] << 118) +
      (src118[60] << 118) +
      (src118[61] << 118) +
      (src118[62] << 118) +
      (src118[63] << 118) +
      (src118[64] << 118) +
      (src118[65] << 118) +
      (src118[66] << 118) +
      (src118[67] << 118) +
      (src118[68] << 118) +
      (src118[69] << 118) +
      (src118[70] << 118) +
      (src118[71] << 118) +
      (src118[72] << 118) +
      (src118[73] << 118) +
      (src118[74] << 118) +
      (src118[75] << 118) +
      (src118[76] << 118) +
      (src118[77] << 118) +
      (src118[78] << 118) +
      (src118[79] << 118) +
      (src118[80] << 118) +
      (src118[81] << 118) +
      (src118[82] << 118) +
      (src118[83] << 118) +
      (src118[84] << 118) +
      (src118[85] << 118) +
      (src118[86] << 118) +
      (src118[87] << 118) +
      (src118[88] << 118) +
      (src118[89] << 118) +
      (src118[90] << 118) +
      (src118[91] << 118) +
      (src118[92] << 118) +
      (src118[93] << 118) +
      (src118[94] << 118) +
      (src118[95] << 118) +
      (src118[96] << 118) +
      (src118[97] << 118) +
      (src118[98] << 118) +
      (src118[99] << 118) +
      (src118[100] << 118) +
      (src118[101] << 118) +
      (src118[102] << 118) +
      (src118[103] << 118) +
      (src118[104] << 118) +
      (src118[105] << 118) +
      (src118[106] << 118) +
      (src118[107] << 118) +
      (src118[108] << 118) +
      (src118[109] << 118) +
      (src118[110] << 118) +
      (src118[111] << 118) +
      (src118[112] << 118) +
      (src118[113] << 118) +
      (src118[114] << 118) +
      (src118[115] << 118) +
      (src118[116] << 118) +
      (src118[117] << 118) +
      (src118[118] << 118) +
      (src118[119] << 118) +
      (src118[120] << 118) +
      (src118[121] << 118) +
      (src118[122] << 118) +
      (src118[123] << 118) +
      (src118[124] << 118) +
      (src118[125] << 118) +
      (src118[126] << 118) +
      (src118[127] << 118) +
      (src119[0] << 119) +
      (src119[1] << 119) +
      (src119[2] << 119) +
      (src119[3] << 119) +
      (src119[4] << 119) +
      (src119[5] << 119) +
      (src119[6] << 119) +
      (src119[7] << 119) +
      (src119[8] << 119) +
      (src119[9] << 119) +
      (src119[10] << 119) +
      (src119[11] << 119) +
      (src119[12] << 119) +
      (src119[13] << 119) +
      (src119[14] << 119) +
      (src119[15] << 119) +
      (src119[16] << 119) +
      (src119[17] << 119) +
      (src119[18] << 119) +
      (src119[19] << 119) +
      (src119[20] << 119) +
      (src119[21] << 119) +
      (src119[22] << 119) +
      (src119[23] << 119) +
      (src119[24] << 119) +
      (src119[25] << 119) +
      (src119[26] << 119) +
      (src119[27] << 119) +
      (src119[28] << 119) +
      (src119[29] << 119) +
      (src119[30] << 119) +
      (src119[31] << 119) +
      (src119[32] << 119) +
      (src119[33] << 119) +
      (src119[34] << 119) +
      (src119[35] << 119) +
      (src119[36] << 119) +
      (src119[37] << 119) +
      (src119[38] << 119) +
      (src119[39] << 119) +
      (src119[40] << 119) +
      (src119[41] << 119) +
      (src119[42] << 119) +
      (src119[43] << 119) +
      (src119[44] << 119) +
      (src119[45] << 119) +
      (src119[46] << 119) +
      (src119[47] << 119) +
      (src119[48] << 119) +
      (src119[49] << 119) +
      (src119[50] << 119) +
      (src119[51] << 119) +
      (src119[52] << 119) +
      (src119[53] << 119) +
      (src119[54] << 119) +
      (src119[55] << 119) +
      (src119[56] << 119) +
      (src119[57] << 119) +
      (src119[58] << 119) +
      (src119[59] << 119) +
      (src119[60] << 119) +
      (src119[61] << 119) +
      (src119[62] << 119) +
      (src119[63] << 119) +
      (src119[64] << 119) +
      (src119[65] << 119) +
      (src119[66] << 119) +
      (src119[67] << 119) +
      (src119[68] << 119) +
      (src119[69] << 119) +
      (src119[70] << 119) +
      (src119[71] << 119) +
      (src119[72] << 119) +
      (src119[73] << 119) +
      (src119[74] << 119) +
      (src119[75] << 119) +
      (src119[76] << 119) +
      (src119[77] << 119) +
      (src119[78] << 119) +
      (src119[79] << 119) +
      (src119[80] << 119) +
      (src119[81] << 119) +
      (src119[82] << 119) +
      (src119[83] << 119) +
      (src119[84] << 119) +
      (src119[85] << 119) +
      (src119[86] << 119) +
      (src119[87] << 119) +
      (src119[88] << 119) +
      (src119[89] << 119) +
      (src119[90] << 119) +
      (src119[91] << 119) +
      (src119[92] << 119) +
      (src119[93] << 119) +
      (src119[94] << 119) +
      (src119[95] << 119) +
      (src119[96] << 119) +
      (src119[97] << 119) +
      (src119[98] << 119) +
      (src119[99] << 119) +
      (src119[100] << 119) +
      (src119[101] << 119) +
      (src119[102] << 119) +
      (src119[103] << 119) +
      (src119[104] << 119) +
      (src119[105] << 119) +
      (src119[106] << 119) +
      (src119[107] << 119) +
      (src119[108] << 119) +
      (src119[109] << 119) +
      (src119[110] << 119) +
      (src119[111] << 119) +
      (src119[112] << 119) +
      (src119[113] << 119) +
      (src119[114] << 119) +
      (src119[115] << 119) +
      (src119[116] << 119) +
      (src119[117] << 119) +
      (src119[118] << 119) +
      (src119[119] << 119) +
      (src119[120] << 119) +
      (src119[121] << 119) +
      (src119[122] << 119) +
      (src119[123] << 119) +
      (src119[124] << 119) +
      (src119[125] << 119) +
      (src119[126] << 119) +
      (src119[127] << 119) +
      (src120[0] << 120) +
      (src120[1] << 120) +
      (src120[2] << 120) +
      (src120[3] << 120) +
      (src120[4] << 120) +
      (src120[5] << 120) +
      (src120[6] << 120) +
      (src120[7] << 120) +
      (src120[8] << 120) +
      (src120[9] << 120) +
      (src120[10] << 120) +
      (src120[11] << 120) +
      (src120[12] << 120) +
      (src120[13] << 120) +
      (src120[14] << 120) +
      (src120[15] << 120) +
      (src120[16] << 120) +
      (src120[17] << 120) +
      (src120[18] << 120) +
      (src120[19] << 120) +
      (src120[20] << 120) +
      (src120[21] << 120) +
      (src120[22] << 120) +
      (src120[23] << 120) +
      (src120[24] << 120) +
      (src120[25] << 120) +
      (src120[26] << 120) +
      (src120[27] << 120) +
      (src120[28] << 120) +
      (src120[29] << 120) +
      (src120[30] << 120) +
      (src120[31] << 120) +
      (src120[32] << 120) +
      (src120[33] << 120) +
      (src120[34] << 120) +
      (src120[35] << 120) +
      (src120[36] << 120) +
      (src120[37] << 120) +
      (src120[38] << 120) +
      (src120[39] << 120) +
      (src120[40] << 120) +
      (src120[41] << 120) +
      (src120[42] << 120) +
      (src120[43] << 120) +
      (src120[44] << 120) +
      (src120[45] << 120) +
      (src120[46] << 120) +
      (src120[47] << 120) +
      (src120[48] << 120) +
      (src120[49] << 120) +
      (src120[50] << 120) +
      (src120[51] << 120) +
      (src120[52] << 120) +
      (src120[53] << 120) +
      (src120[54] << 120) +
      (src120[55] << 120) +
      (src120[56] << 120) +
      (src120[57] << 120) +
      (src120[58] << 120) +
      (src120[59] << 120) +
      (src120[60] << 120) +
      (src120[61] << 120) +
      (src120[62] << 120) +
      (src120[63] << 120) +
      (src120[64] << 120) +
      (src120[65] << 120) +
      (src120[66] << 120) +
      (src120[67] << 120) +
      (src120[68] << 120) +
      (src120[69] << 120) +
      (src120[70] << 120) +
      (src120[71] << 120) +
      (src120[72] << 120) +
      (src120[73] << 120) +
      (src120[74] << 120) +
      (src120[75] << 120) +
      (src120[76] << 120) +
      (src120[77] << 120) +
      (src120[78] << 120) +
      (src120[79] << 120) +
      (src120[80] << 120) +
      (src120[81] << 120) +
      (src120[82] << 120) +
      (src120[83] << 120) +
      (src120[84] << 120) +
      (src120[85] << 120) +
      (src120[86] << 120) +
      (src120[87] << 120) +
      (src120[88] << 120) +
      (src120[89] << 120) +
      (src120[90] << 120) +
      (src120[91] << 120) +
      (src120[92] << 120) +
      (src120[93] << 120) +
      (src120[94] << 120) +
      (src120[95] << 120) +
      (src120[96] << 120) +
      (src120[97] << 120) +
      (src120[98] << 120) +
      (src120[99] << 120) +
      (src120[100] << 120) +
      (src120[101] << 120) +
      (src120[102] << 120) +
      (src120[103] << 120) +
      (src120[104] << 120) +
      (src120[105] << 120) +
      (src120[106] << 120) +
      (src120[107] << 120) +
      (src120[108] << 120) +
      (src120[109] << 120) +
      (src120[110] << 120) +
      (src120[111] << 120) +
      (src120[112] << 120) +
      (src120[113] << 120) +
      (src120[114] << 120) +
      (src120[115] << 120) +
      (src120[116] << 120) +
      (src120[117] << 120) +
      (src120[118] << 120) +
      (src120[119] << 120) +
      (src120[120] << 120) +
      (src120[121] << 120) +
      (src120[122] << 120) +
      (src120[123] << 120) +
      (src120[124] << 120) +
      (src120[125] << 120) +
      (src120[126] << 120) +
      (src120[127] << 120) +
      (src121[0] << 121) +
      (src121[1] << 121) +
      (src121[2] << 121) +
      (src121[3] << 121) +
      (src121[4] << 121) +
      (src121[5] << 121) +
      (src121[6] << 121) +
      (src121[7] << 121) +
      (src121[8] << 121) +
      (src121[9] << 121) +
      (src121[10] << 121) +
      (src121[11] << 121) +
      (src121[12] << 121) +
      (src121[13] << 121) +
      (src121[14] << 121) +
      (src121[15] << 121) +
      (src121[16] << 121) +
      (src121[17] << 121) +
      (src121[18] << 121) +
      (src121[19] << 121) +
      (src121[20] << 121) +
      (src121[21] << 121) +
      (src121[22] << 121) +
      (src121[23] << 121) +
      (src121[24] << 121) +
      (src121[25] << 121) +
      (src121[26] << 121) +
      (src121[27] << 121) +
      (src121[28] << 121) +
      (src121[29] << 121) +
      (src121[30] << 121) +
      (src121[31] << 121) +
      (src121[32] << 121) +
      (src121[33] << 121) +
      (src121[34] << 121) +
      (src121[35] << 121) +
      (src121[36] << 121) +
      (src121[37] << 121) +
      (src121[38] << 121) +
      (src121[39] << 121) +
      (src121[40] << 121) +
      (src121[41] << 121) +
      (src121[42] << 121) +
      (src121[43] << 121) +
      (src121[44] << 121) +
      (src121[45] << 121) +
      (src121[46] << 121) +
      (src121[47] << 121) +
      (src121[48] << 121) +
      (src121[49] << 121) +
      (src121[50] << 121) +
      (src121[51] << 121) +
      (src121[52] << 121) +
      (src121[53] << 121) +
      (src121[54] << 121) +
      (src121[55] << 121) +
      (src121[56] << 121) +
      (src121[57] << 121) +
      (src121[58] << 121) +
      (src121[59] << 121) +
      (src121[60] << 121) +
      (src121[61] << 121) +
      (src121[62] << 121) +
      (src121[63] << 121) +
      (src121[64] << 121) +
      (src121[65] << 121) +
      (src121[66] << 121) +
      (src121[67] << 121) +
      (src121[68] << 121) +
      (src121[69] << 121) +
      (src121[70] << 121) +
      (src121[71] << 121) +
      (src121[72] << 121) +
      (src121[73] << 121) +
      (src121[74] << 121) +
      (src121[75] << 121) +
      (src121[76] << 121) +
      (src121[77] << 121) +
      (src121[78] << 121) +
      (src121[79] << 121) +
      (src121[80] << 121) +
      (src121[81] << 121) +
      (src121[82] << 121) +
      (src121[83] << 121) +
      (src121[84] << 121) +
      (src121[85] << 121) +
      (src121[86] << 121) +
      (src121[87] << 121) +
      (src121[88] << 121) +
      (src121[89] << 121) +
      (src121[90] << 121) +
      (src121[91] << 121) +
      (src121[92] << 121) +
      (src121[93] << 121) +
      (src121[94] << 121) +
      (src121[95] << 121) +
      (src121[96] << 121) +
      (src121[97] << 121) +
      (src121[98] << 121) +
      (src121[99] << 121) +
      (src121[100] << 121) +
      (src121[101] << 121) +
      (src121[102] << 121) +
      (src121[103] << 121) +
      (src121[104] << 121) +
      (src121[105] << 121) +
      (src121[106] << 121) +
      (src121[107] << 121) +
      (src121[108] << 121) +
      (src121[109] << 121) +
      (src121[110] << 121) +
      (src121[111] << 121) +
      (src121[112] << 121) +
      (src121[113] << 121) +
      (src121[114] << 121) +
      (src121[115] << 121) +
      (src121[116] << 121) +
      (src121[117] << 121) +
      (src121[118] << 121) +
      (src121[119] << 121) +
      (src121[120] << 121) +
      (src121[121] << 121) +
      (src121[122] << 121) +
      (src121[123] << 121) +
      (src121[124] << 121) +
      (src121[125] << 121) +
      (src121[126] << 121) +
      (src121[127] << 121) +
      (src122[0] << 122) +
      (src122[1] << 122) +
      (src122[2] << 122) +
      (src122[3] << 122) +
      (src122[4] << 122) +
      (src122[5] << 122) +
      (src122[6] << 122) +
      (src122[7] << 122) +
      (src122[8] << 122) +
      (src122[9] << 122) +
      (src122[10] << 122) +
      (src122[11] << 122) +
      (src122[12] << 122) +
      (src122[13] << 122) +
      (src122[14] << 122) +
      (src122[15] << 122) +
      (src122[16] << 122) +
      (src122[17] << 122) +
      (src122[18] << 122) +
      (src122[19] << 122) +
      (src122[20] << 122) +
      (src122[21] << 122) +
      (src122[22] << 122) +
      (src122[23] << 122) +
      (src122[24] << 122) +
      (src122[25] << 122) +
      (src122[26] << 122) +
      (src122[27] << 122) +
      (src122[28] << 122) +
      (src122[29] << 122) +
      (src122[30] << 122) +
      (src122[31] << 122) +
      (src122[32] << 122) +
      (src122[33] << 122) +
      (src122[34] << 122) +
      (src122[35] << 122) +
      (src122[36] << 122) +
      (src122[37] << 122) +
      (src122[38] << 122) +
      (src122[39] << 122) +
      (src122[40] << 122) +
      (src122[41] << 122) +
      (src122[42] << 122) +
      (src122[43] << 122) +
      (src122[44] << 122) +
      (src122[45] << 122) +
      (src122[46] << 122) +
      (src122[47] << 122) +
      (src122[48] << 122) +
      (src122[49] << 122) +
      (src122[50] << 122) +
      (src122[51] << 122) +
      (src122[52] << 122) +
      (src122[53] << 122) +
      (src122[54] << 122) +
      (src122[55] << 122) +
      (src122[56] << 122) +
      (src122[57] << 122) +
      (src122[58] << 122) +
      (src122[59] << 122) +
      (src122[60] << 122) +
      (src122[61] << 122) +
      (src122[62] << 122) +
      (src122[63] << 122) +
      (src122[64] << 122) +
      (src122[65] << 122) +
      (src122[66] << 122) +
      (src122[67] << 122) +
      (src122[68] << 122) +
      (src122[69] << 122) +
      (src122[70] << 122) +
      (src122[71] << 122) +
      (src122[72] << 122) +
      (src122[73] << 122) +
      (src122[74] << 122) +
      (src122[75] << 122) +
      (src122[76] << 122) +
      (src122[77] << 122) +
      (src122[78] << 122) +
      (src122[79] << 122) +
      (src122[80] << 122) +
      (src122[81] << 122) +
      (src122[82] << 122) +
      (src122[83] << 122) +
      (src122[84] << 122) +
      (src122[85] << 122) +
      (src122[86] << 122) +
      (src122[87] << 122) +
      (src122[88] << 122) +
      (src122[89] << 122) +
      (src122[90] << 122) +
      (src122[91] << 122) +
      (src122[92] << 122) +
      (src122[93] << 122) +
      (src122[94] << 122) +
      (src122[95] << 122) +
      (src122[96] << 122) +
      (src122[97] << 122) +
      (src122[98] << 122) +
      (src122[99] << 122) +
      (src122[100] << 122) +
      (src122[101] << 122) +
      (src122[102] << 122) +
      (src122[103] << 122) +
      (src122[104] << 122) +
      (src122[105] << 122) +
      (src122[106] << 122) +
      (src122[107] << 122) +
      (src122[108] << 122) +
      (src122[109] << 122) +
      (src122[110] << 122) +
      (src122[111] << 122) +
      (src122[112] << 122) +
      (src122[113] << 122) +
      (src122[114] << 122) +
      (src122[115] << 122) +
      (src122[116] << 122) +
      (src122[117] << 122) +
      (src122[118] << 122) +
      (src122[119] << 122) +
      (src122[120] << 122) +
      (src122[121] << 122) +
      (src122[122] << 122) +
      (src122[123] << 122) +
      (src122[124] << 122) +
      (src122[125] << 122) +
      (src122[126] << 122) +
      (src122[127] << 122) +
      (src123[0] << 123) +
      (src123[1] << 123) +
      (src123[2] << 123) +
      (src123[3] << 123) +
      (src123[4] << 123) +
      (src123[5] << 123) +
      (src123[6] << 123) +
      (src123[7] << 123) +
      (src123[8] << 123) +
      (src123[9] << 123) +
      (src123[10] << 123) +
      (src123[11] << 123) +
      (src123[12] << 123) +
      (src123[13] << 123) +
      (src123[14] << 123) +
      (src123[15] << 123) +
      (src123[16] << 123) +
      (src123[17] << 123) +
      (src123[18] << 123) +
      (src123[19] << 123) +
      (src123[20] << 123) +
      (src123[21] << 123) +
      (src123[22] << 123) +
      (src123[23] << 123) +
      (src123[24] << 123) +
      (src123[25] << 123) +
      (src123[26] << 123) +
      (src123[27] << 123) +
      (src123[28] << 123) +
      (src123[29] << 123) +
      (src123[30] << 123) +
      (src123[31] << 123) +
      (src123[32] << 123) +
      (src123[33] << 123) +
      (src123[34] << 123) +
      (src123[35] << 123) +
      (src123[36] << 123) +
      (src123[37] << 123) +
      (src123[38] << 123) +
      (src123[39] << 123) +
      (src123[40] << 123) +
      (src123[41] << 123) +
      (src123[42] << 123) +
      (src123[43] << 123) +
      (src123[44] << 123) +
      (src123[45] << 123) +
      (src123[46] << 123) +
      (src123[47] << 123) +
      (src123[48] << 123) +
      (src123[49] << 123) +
      (src123[50] << 123) +
      (src123[51] << 123) +
      (src123[52] << 123) +
      (src123[53] << 123) +
      (src123[54] << 123) +
      (src123[55] << 123) +
      (src123[56] << 123) +
      (src123[57] << 123) +
      (src123[58] << 123) +
      (src123[59] << 123) +
      (src123[60] << 123) +
      (src123[61] << 123) +
      (src123[62] << 123) +
      (src123[63] << 123) +
      (src123[64] << 123) +
      (src123[65] << 123) +
      (src123[66] << 123) +
      (src123[67] << 123) +
      (src123[68] << 123) +
      (src123[69] << 123) +
      (src123[70] << 123) +
      (src123[71] << 123) +
      (src123[72] << 123) +
      (src123[73] << 123) +
      (src123[74] << 123) +
      (src123[75] << 123) +
      (src123[76] << 123) +
      (src123[77] << 123) +
      (src123[78] << 123) +
      (src123[79] << 123) +
      (src123[80] << 123) +
      (src123[81] << 123) +
      (src123[82] << 123) +
      (src123[83] << 123) +
      (src123[84] << 123) +
      (src123[85] << 123) +
      (src123[86] << 123) +
      (src123[87] << 123) +
      (src123[88] << 123) +
      (src123[89] << 123) +
      (src123[90] << 123) +
      (src123[91] << 123) +
      (src123[92] << 123) +
      (src123[93] << 123) +
      (src123[94] << 123) +
      (src123[95] << 123) +
      (src123[96] << 123) +
      (src123[97] << 123) +
      (src123[98] << 123) +
      (src123[99] << 123) +
      (src123[100] << 123) +
      (src123[101] << 123) +
      (src123[102] << 123) +
      (src123[103] << 123) +
      (src123[104] << 123) +
      (src123[105] << 123) +
      (src123[106] << 123) +
      (src123[107] << 123) +
      (src123[108] << 123) +
      (src123[109] << 123) +
      (src123[110] << 123) +
      (src123[111] << 123) +
      (src123[112] << 123) +
      (src123[113] << 123) +
      (src123[114] << 123) +
      (src123[115] << 123) +
      (src123[116] << 123) +
      (src123[117] << 123) +
      (src123[118] << 123) +
      (src123[119] << 123) +
      (src123[120] << 123) +
      (src123[121] << 123) +
      (src123[122] << 123) +
      (src123[123] << 123) +
      (src123[124] << 123) +
      (src123[125] << 123) +
      (src123[126] << 123) +
      (src123[127] << 123) +
      (src124[0] << 124) +
      (src124[1] << 124) +
      (src124[2] << 124) +
      (src124[3] << 124) +
      (src124[4] << 124) +
      (src124[5] << 124) +
      (src124[6] << 124) +
      (src124[7] << 124) +
      (src124[8] << 124) +
      (src124[9] << 124) +
      (src124[10] << 124) +
      (src124[11] << 124) +
      (src124[12] << 124) +
      (src124[13] << 124) +
      (src124[14] << 124) +
      (src124[15] << 124) +
      (src124[16] << 124) +
      (src124[17] << 124) +
      (src124[18] << 124) +
      (src124[19] << 124) +
      (src124[20] << 124) +
      (src124[21] << 124) +
      (src124[22] << 124) +
      (src124[23] << 124) +
      (src124[24] << 124) +
      (src124[25] << 124) +
      (src124[26] << 124) +
      (src124[27] << 124) +
      (src124[28] << 124) +
      (src124[29] << 124) +
      (src124[30] << 124) +
      (src124[31] << 124) +
      (src124[32] << 124) +
      (src124[33] << 124) +
      (src124[34] << 124) +
      (src124[35] << 124) +
      (src124[36] << 124) +
      (src124[37] << 124) +
      (src124[38] << 124) +
      (src124[39] << 124) +
      (src124[40] << 124) +
      (src124[41] << 124) +
      (src124[42] << 124) +
      (src124[43] << 124) +
      (src124[44] << 124) +
      (src124[45] << 124) +
      (src124[46] << 124) +
      (src124[47] << 124) +
      (src124[48] << 124) +
      (src124[49] << 124) +
      (src124[50] << 124) +
      (src124[51] << 124) +
      (src124[52] << 124) +
      (src124[53] << 124) +
      (src124[54] << 124) +
      (src124[55] << 124) +
      (src124[56] << 124) +
      (src124[57] << 124) +
      (src124[58] << 124) +
      (src124[59] << 124) +
      (src124[60] << 124) +
      (src124[61] << 124) +
      (src124[62] << 124) +
      (src124[63] << 124) +
      (src124[64] << 124) +
      (src124[65] << 124) +
      (src124[66] << 124) +
      (src124[67] << 124) +
      (src124[68] << 124) +
      (src124[69] << 124) +
      (src124[70] << 124) +
      (src124[71] << 124) +
      (src124[72] << 124) +
      (src124[73] << 124) +
      (src124[74] << 124) +
      (src124[75] << 124) +
      (src124[76] << 124) +
      (src124[77] << 124) +
      (src124[78] << 124) +
      (src124[79] << 124) +
      (src124[80] << 124) +
      (src124[81] << 124) +
      (src124[82] << 124) +
      (src124[83] << 124) +
      (src124[84] << 124) +
      (src124[85] << 124) +
      (src124[86] << 124) +
      (src124[87] << 124) +
      (src124[88] << 124) +
      (src124[89] << 124) +
      (src124[90] << 124) +
      (src124[91] << 124) +
      (src124[92] << 124) +
      (src124[93] << 124) +
      (src124[94] << 124) +
      (src124[95] << 124) +
      (src124[96] << 124) +
      (src124[97] << 124) +
      (src124[98] << 124) +
      (src124[99] << 124) +
      (src124[100] << 124) +
      (src124[101] << 124) +
      (src124[102] << 124) +
      (src124[103] << 124) +
      (src124[104] << 124) +
      (src124[105] << 124) +
      (src124[106] << 124) +
      (src124[107] << 124) +
      (src124[108] << 124) +
      (src124[109] << 124) +
      (src124[110] << 124) +
      (src124[111] << 124) +
      (src124[112] << 124) +
      (src124[113] << 124) +
      (src124[114] << 124) +
      (src124[115] << 124) +
      (src124[116] << 124) +
      (src124[117] << 124) +
      (src124[118] << 124) +
      (src124[119] << 124) +
      (src124[120] << 124) +
      (src124[121] << 124) +
      (src124[122] << 124) +
      (src124[123] << 124) +
      (src124[124] << 124) +
      (src124[125] << 124) +
      (src124[126] << 124) +
      (src124[127] << 124) +
      (src125[0] << 125) +
      (src125[1] << 125) +
      (src125[2] << 125) +
      (src125[3] << 125) +
      (src125[4] << 125) +
      (src125[5] << 125) +
      (src125[6] << 125) +
      (src125[7] << 125) +
      (src125[8] << 125) +
      (src125[9] << 125) +
      (src125[10] << 125) +
      (src125[11] << 125) +
      (src125[12] << 125) +
      (src125[13] << 125) +
      (src125[14] << 125) +
      (src125[15] << 125) +
      (src125[16] << 125) +
      (src125[17] << 125) +
      (src125[18] << 125) +
      (src125[19] << 125) +
      (src125[20] << 125) +
      (src125[21] << 125) +
      (src125[22] << 125) +
      (src125[23] << 125) +
      (src125[24] << 125) +
      (src125[25] << 125) +
      (src125[26] << 125) +
      (src125[27] << 125) +
      (src125[28] << 125) +
      (src125[29] << 125) +
      (src125[30] << 125) +
      (src125[31] << 125) +
      (src125[32] << 125) +
      (src125[33] << 125) +
      (src125[34] << 125) +
      (src125[35] << 125) +
      (src125[36] << 125) +
      (src125[37] << 125) +
      (src125[38] << 125) +
      (src125[39] << 125) +
      (src125[40] << 125) +
      (src125[41] << 125) +
      (src125[42] << 125) +
      (src125[43] << 125) +
      (src125[44] << 125) +
      (src125[45] << 125) +
      (src125[46] << 125) +
      (src125[47] << 125) +
      (src125[48] << 125) +
      (src125[49] << 125) +
      (src125[50] << 125) +
      (src125[51] << 125) +
      (src125[52] << 125) +
      (src125[53] << 125) +
      (src125[54] << 125) +
      (src125[55] << 125) +
      (src125[56] << 125) +
      (src125[57] << 125) +
      (src125[58] << 125) +
      (src125[59] << 125) +
      (src125[60] << 125) +
      (src125[61] << 125) +
      (src125[62] << 125) +
      (src125[63] << 125) +
      (src125[64] << 125) +
      (src125[65] << 125) +
      (src125[66] << 125) +
      (src125[67] << 125) +
      (src125[68] << 125) +
      (src125[69] << 125) +
      (src125[70] << 125) +
      (src125[71] << 125) +
      (src125[72] << 125) +
      (src125[73] << 125) +
      (src125[74] << 125) +
      (src125[75] << 125) +
      (src125[76] << 125) +
      (src125[77] << 125) +
      (src125[78] << 125) +
      (src125[79] << 125) +
      (src125[80] << 125) +
      (src125[81] << 125) +
      (src125[82] << 125) +
      (src125[83] << 125) +
      (src125[84] << 125) +
      (src125[85] << 125) +
      (src125[86] << 125) +
      (src125[87] << 125) +
      (src125[88] << 125) +
      (src125[89] << 125) +
      (src125[90] << 125) +
      (src125[91] << 125) +
      (src125[92] << 125) +
      (src125[93] << 125) +
      (src125[94] << 125) +
      (src125[95] << 125) +
      (src125[96] << 125) +
      (src125[97] << 125) +
      (src125[98] << 125) +
      (src125[99] << 125) +
      (src125[100] << 125) +
      (src125[101] << 125) +
      (src125[102] << 125) +
      (src125[103] << 125) +
      (src125[104] << 125) +
      (src125[105] << 125) +
      (src125[106] << 125) +
      (src125[107] << 125) +
      (src125[108] << 125) +
      (src125[109] << 125) +
      (src125[110] << 125) +
      (src125[111] << 125) +
      (src125[112] << 125) +
      (src125[113] << 125) +
      (src125[114] << 125) +
      (src125[115] << 125) +
      (src125[116] << 125) +
      (src125[117] << 125) +
      (src125[118] << 125) +
      (src125[119] << 125) +
      (src125[120] << 125) +
      (src125[121] << 125) +
      (src125[122] << 125) +
      (src125[123] << 125) +
      (src125[124] << 125) +
      (src125[125] << 125) +
      (src125[126] << 125) +
      (src125[127] << 125) +
      (src126[0] << 126) +
      (src126[1] << 126) +
      (src126[2] << 126) +
      (src126[3] << 126) +
      (src126[4] << 126) +
      (src126[5] << 126) +
      (src126[6] << 126) +
      (src126[7] << 126) +
      (src126[8] << 126) +
      (src126[9] << 126) +
      (src126[10] << 126) +
      (src126[11] << 126) +
      (src126[12] << 126) +
      (src126[13] << 126) +
      (src126[14] << 126) +
      (src126[15] << 126) +
      (src126[16] << 126) +
      (src126[17] << 126) +
      (src126[18] << 126) +
      (src126[19] << 126) +
      (src126[20] << 126) +
      (src126[21] << 126) +
      (src126[22] << 126) +
      (src126[23] << 126) +
      (src126[24] << 126) +
      (src126[25] << 126) +
      (src126[26] << 126) +
      (src126[27] << 126) +
      (src126[28] << 126) +
      (src126[29] << 126) +
      (src126[30] << 126) +
      (src126[31] << 126) +
      (src126[32] << 126) +
      (src126[33] << 126) +
      (src126[34] << 126) +
      (src126[35] << 126) +
      (src126[36] << 126) +
      (src126[37] << 126) +
      (src126[38] << 126) +
      (src126[39] << 126) +
      (src126[40] << 126) +
      (src126[41] << 126) +
      (src126[42] << 126) +
      (src126[43] << 126) +
      (src126[44] << 126) +
      (src126[45] << 126) +
      (src126[46] << 126) +
      (src126[47] << 126) +
      (src126[48] << 126) +
      (src126[49] << 126) +
      (src126[50] << 126) +
      (src126[51] << 126) +
      (src126[52] << 126) +
      (src126[53] << 126) +
      (src126[54] << 126) +
      (src126[55] << 126) +
      (src126[56] << 126) +
      (src126[57] << 126) +
      (src126[58] << 126) +
      (src126[59] << 126) +
      (src126[60] << 126) +
      (src126[61] << 126) +
      (src126[62] << 126) +
      (src126[63] << 126) +
      (src126[64] << 126) +
      (src126[65] << 126) +
      (src126[66] << 126) +
      (src126[67] << 126) +
      (src126[68] << 126) +
      (src126[69] << 126) +
      (src126[70] << 126) +
      (src126[71] << 126) +
      (src126[72] << 126) +
      (src126[73] << 126) +
      (src126[74] << 126) +
      (src126[75] << 126) +
      (src126[76] << 126) +
      (src126[77] << 126) +
      (src126[78] << 126) +
      (src126[79] << 126) +
      (src126[80] << 126) +
      (src126[81] << 126) +
      (src126[82] << 126) +
      (src126[83] << 126) +
      (src126[84] << 126) +
      (src126[85] << 126) +
      (src126[86] << 126) +
      (src126[87] << 126) +
      (src126[88] << 126) +
      (src126[89] << 126) +
      (src126[90] << 126) +
      (src126[91] << 126) +
      (src126[92] << 126) +
      (src126[93] << 126) +
      (src126[94] << 126) +
      (src126[95] << 126) +
      (src126[96] << 126) +
      (src126[97] << 126) +
      (src126[98] << 126) +
      (src126[99] << 126) +
      (src126[100] << 126) +
      (src126[101] << 126) +
      (src126[102] << 126) +
      (src126[103] << 126) +
      (src126[104] << 126) +
      (src126[105] << 126) +
      (src126[106] << 126) +
      (src126[107] << 126) +
      (src126[108] << 126) +
      (src126[109] << 126) +
      (src126[110] << 126) +
      (src126[111] << 126) +
      (src126[112] << 126) +
      (src126[113] << 126) +
      (src126[114] << 126) +
      (src126[115] << 126) +
      (src126[116] << 126) +
      (src126[117] << 126) +
      (src126[118] << 126) +
      (src126[119] << 126) +
      (src126[120] << 126) +
      (src126[121] << 126) +
      (src126[122] << 126) +
      (src126[123] << 126) +
      (src126[124] << 126) +
      (src126[125] << 126) +
      (src126[126] << 126) +
      (src126[127] << 126) +
      (src127[0] << 127) +
      (src127[1] << 127) +
      (src127[2] << 127) +
      (src127[3] << 127) +
      (src127[4] << 127) +
      (src127[5] << 127) +
      (src127[6] << 127) +
      (src127[7] << 127) +
      (src127[8] << 127) +
      (src127[9] << 127) +
      (src127[10] << 127) +
      (src127[11] << 127) +
      (src127[12] << 127) +
      (src127[13] << 127) +
      (src127[14] << 127) +
      (src127[15] << 127) +
      (src127[16] << 127) +
      (src127[17] << 127) +
      (src127[18] << 127) +
      (src127[19] << 127) +
      (src127[20] << 127) +
      (src127[21] << 127) +
      (src127[22] << 127) +
      (src127[23] << 127) +
      (src127[24] << 127) +
      (src127[25] << 127) +
      (src127[26] << 127) +
      (src127[27] << 127) +
      (src127[28] << 127) +
      (src127[29] << 127) +
      (src127[30] << 127) +
      (src127[31] << 127) +
      (src127[32] << 127) +
      (src127[33] << 127) +
      (src127[34] << 127) +
      (src127[35] << 127) +
      (src127[36] << 127) +
      (src127[37] << 127) +
      (src127[38] << 127) +
      (src127[39] << 127) +
      (src127[40] << 127) +
      (src127[41] << 127) +
      (src127[42] << 127) +
      (src127[43] << 127) +
      (src127[44] << 127) +
      (src127[45] << 127) +
      (src127[46] << 127) +
      (src127[47] << 127) +
      (src127[48] << 127) +
      (src127[49] << 127) +
      (src127[50] << 127) +
      (src127[51] << 127) +
      (src127[52] << 127) +
      (src127[53] << 127) +
      (src127[54] << 127) +
      (src127[55] << 127) +
      (src127[56] << 127) +
      (src127[57] << 127) +
      (src127[58] << 127) +
      (src127[59] << 127) +
      (src127[60] << 127) +
      (src127[61] << 127) +
      (src127[62] << 127) +
      (src127[63] << 127) +
      (src127[64] << 127) +
      (src127[65] << 127) +
      (src127[66] << 127) +
      (src127[67] << 127) +
      (src127[68] << 127) +
      (src127[69] << 127) +
      (src127[70] << 127) +
      (src127[71] << 127) +
      (src127[72] << 127) +
      (src127[73] << 127) +
      (src127[74] << 127) +
      (src127[75] << 127) +
      (src127[76] << 127) +
      (src127[77] << 127) +
      (src127[78] << 127) +
      (src127[79] << 127) +
      (src127[80] << 127) +
      (src127[81] << 127) +
      (src127[82] << 127) +
      (src127[83] << 127) +
      (src127[84] << 127) +
      (src127[85] << 127) +
      (src127[86] << 127) +
      (src127[87] << 127) +
      (src127[88] << 127) +
      (src127[89] << 127) +
      (src127[90] << 127) +
      (src127[91] << 127) +
      (src127[92] << 127) +
      (src127[93] << 127) +
      (src127[94] << 127) +
      (src127[95] << 127) +
      (src127[96] << 127) +
      (src127[97] << 127) +
      (src127[98] << 127) +
      (src127[99] << 127) +
      (src127[100] << 127) +
      (src127[101] << 127) +
      (src127[102] << 127) +
      (src127[103] << 127) +
      (src127[104] << 127) +
      (src127[105] << 127) +
      (src127[106] << 127) +
      (src127[107] << 127) +
      (src127[108] << 127) +
      (src127[109] << 127) +
      (src127[110] << 127) +
      (src127[111] << 127) +
      (src127[112] << 127) +
      (src127[113] << 127) +
      (src127[114] << 127) +
      (src127[115] << 127) +
      (src127[116] << 127) +
      (src127[117] << 127) +
      (src127[118] << 127) +
      (src127[119] << 127) +
      (src127[120] << 127) +
      (src127[121] << 127) +
      (src127[122] << 127) +
      (src127[123] << 127) +
      (src127[124] << 127) +
      (src127[125] << 127) +
      (src127[126] << 127) +
      (src127[127] << 127);
   assign dstsum =
      (dst000[0] << 0) +
      (dst000[1] << 0) +
      (dst001[0] << 1) +
      (dst001[1] << 1) +
      (dst002[0] << 2) +
      (dst002[1] << 2) +
      (dst003[0] << 3) +
      (dst004[0] << 4) +
      (dst005[0] << 5) +
      (dst005[1] << 5) +
      (dst006[0] << 6) +
      (dst007[0] << 7) +
      (dst007[1] << 7) +
      (dst008[0] << 8) +
      (dst008[1] << 8) +
      (dst009[0] << 9) +
      (dst009[1] << 9) +
      (dst010[0] << 10) +
      (dst010[1] << 10) +
      (dst011[0] << 11) +
      (dst011[1] << 11) +
      (dst012[0] << 12) +
      (dst012[1] << 12) +
      (dst013[0] << 13) +
      (dst014[0] << 14) +
      (dst014[1] << 14) +
      (dst015[0] << 15) +
      (dst015[1] << 15) +
      (dst016[0] << 16) +
      (dst016[1] << 16) +
      (dst017[0] << 17) +
      (dst017[1] << 17) +
      (dst018[0] << 18) +
      (dst018[1] << 18) +
      (dst019[0] << 19) +
      (dst019[1] << 19) +
      (dst020[0] << 20) +
      (dst020[1] << 20) +
      (dst021[0] << 21) +
      (dst021[1] << 21) +
      (dst022[0] << 22) +
      (dst022[1] << 22) +
      (dst023[0] << 23) +
      (dst023[1] << 23) +
      (dst024[0] << 24) +
      (dst024[1] << 24) +
      (dst025[0] << 25) +
      (dst025[1] << 25) +
      (dst026[0] << 26) +
      (dst026[1] << 26) +
      (dst027[0] << 27) +
      (dst027[1] << 27) +
      (dst028[0] << 28) +
      (dst028[1] << 28) +
      (dst029[0] << 29) +
      (dst029[1] << 29) +
      (dst030[0] << 30) +
      (dst030[1] << 30) +
      (dst031[0] << 31) +
      (dst031[1] << 31) +
      (dst032[0] << 32) +
      (dst032[1] << 32) +
      (dst033[0] << 33) +
      (dst033[1] << 33) +
      (dst034[0] << 34) +
      (dst034[1] << 34) +
      (dst035[0] << 35) +
      (dst035[1] << 35) +
      (dst036[0] << 36) +
      (dst036[1] << 36) +
      (dst037[0] << 37) +
      (dst037[1] << 37) +
      (dst038[0] << 38) +
      (dst039[0] << 39) +
      (dst040[0] << 40) +
      (dst040[1] << 40) +
      (dst041[0] << 41) +
      (dst041[1] << 41) +
      (dst042[0] << 42) +
      (dst042[1] << 42) +
      (dst043[0] << 43) +
      (dst043[1] << 43) +
      (dst044[0] << 44) +
      (dst044[1] << 44) +
      (dst045[0] << 45) +
      (dst045[1] << 45) +
      (dst046[0] << 46) +
      (dst046[1] << 46) +
      (dst047[0] << 47) +
      (dst047[1] << 47) +
      (dst048[0] << 48) +
      (dst048[1] << 48) +
      (dst049[0] << 49) +
      (dst049[1] << 49) +
      (dst050[0] << 50) +
      (dst050[1] << 50) +
      (dst051[0] << 51) +
      (dst051[1] << 51) +
      (dst052[0] << 52) +
      (dst052[1] << 52) +
      (dst053[0] << 53) +
      (dst053[1] << 53) +
      (dst054[0] << 54) +
      (dst054[1] << 54) +
      (dst055[0] << 55) +
      (dst055[1] << 55) +
      (dst056[0] << 56) +
      (dst056[1] << 56) +
      (dst057[0] << 57) +
      (dst057[1] << 57) +
      (dst058[0] << 58) +
      (dst058[1] << 58) +
      (dst059[0] << 59) +
      (dst059[1] << 59) +
      (dst060[0] << 60) +
      (dst060[1] << 60) +
      (dst061[0] << 61) +
      (dst062[0] << 62) +
      (dst062[1] << 62) +
      (dst063[0] << 63) +
      (dst063[1] << 63) +
      (dst064[0] << 64) +
      (dst064[1] << 64) +
      (dst065[0] << 65) +
      (dst065[1] << 65) +
      (dst066[0] << 66) +
      (dst066[1] << 66) +
      (dst067[0] << 67) +
      (dst068[0] << 68) +
      (dst068[1] << 68) +
      (dst069[0] << 69) +
      (dst069[1] << 69) +
      (dst070[0] << 70) +
      (dst070[1] << 70) +
      (dst071[0] << 71) +
      (dst071[1] << 71) +
      (dst072[0] << 72) +
      (dst072[1] << 72) +
      (dst073[0] << 73) +
      (dst073[1] << 73) +
      (dst074[0] << 74) +
      (dst074[1] << 74) +
      (dst075[0] << 75) +
      (dst075[1] << 75) +
      (dst076[0] << 76) +
      (dst076[1] << 76) +
      (dst077[0] << 77) +
      (dst077[1] << 77) +
      (dst078[0] << 78) +
      (dst078[1] << 78) +
      (dst079[0] << 79) +
      (dst079[1] << 79) +
      (dst080[0] << 80) +
      (dst080[1] << 80) +
      (dst081[0] << 81) +
      (dst081[1] << 81) +
      (dst082[0] << 82) +
      (dst082[1] << 82) +
      (dst083[0] << 83) +
      (dst084[0] << 84) +
      (dst084[1] << 84) +
      (dst085[0] << 85) +
      (dst085[1] << 85) +
      (dst086[0] << 86) +
      (dst086[1] << 86) +
      (dst087[0] << 87) +
      (dst087[1] << 87) +
      (dst088[0] << 88) +
      (dst088[1] << 88) +
      (dst089[0] << 89) +
      (dst089[1] << 89) +
      (dst090[0] << 90) +
      (dst090[1] << 90) +
      (dst091[0] << 91) +
      (dst091[1] << 91) +
      (dst092[0] << 92) +
      (dst092[1] << 92) +
      (dst093[0] << 93) +
      (dst093[1] << 93) +
      (dst094[0] << 94) +
      (dst094[1] << 94) +
      (dst095[0] << 95) +
      (dst095[1] << 95) +
      (dst096[0] << 96) +
      (dst096[1] << 96) +
      (dst097[0] << 97) +
      (dst097[1] << 97) +
      (dst098[0] << 98) +
      (dst098[1] << 98) +
      (dst099[0] << 99) +
      (dst099[1] << 99) +
      (dst100[0] << 100) +
      (dst100[1] << 100) +
      (dst101[0] << 101) +
      (dst101[1] << 101) +
      (dst102[0] << 102) +
      (dst102[1] << 102) +
      (dst103[0] << 103) +
      (dst103[1] << 103) +
      (dst104[0] << 104) +
      (dst104[1] << 104) +
      (dst105[0] << 105) +
      (dst105[1] << 105) +
      (dst106[0] << 106) +
      (dst106[1] << 106) +
      (dst107[0] << 107) +
      (dst107[1] << 107) +
      (dst108[0] << 108) +
      (dst108[1] << 108) +
      (dst109[0] << 109) +
      (dst109[1] << 109) +
      (dst110[0] << 110) +
      (dst110[1] << 110) +
      (dst111[0] << 111) +
      (dst111[1] << 111) +
      (dst112[0] << 112) +
      (dst113[0] << 113) +
      (dst113[1] << 113) +
      (dst114[0] << 114) +
      (dst114[1] << 114) +
      (dst115[0] << 115) +
      (dst115[1] << 115) +
      (dst116[0] << 116) +
      (dst116[1] << 116) +
      (dst117[0] << 117) +
      (dst117[1] << 117) +
      (dst118[0] << 118) +
      (dst118[1] << 118) +
      (dst119[0] << 119) +
      (dst119[1] << 119) +
      (dst120[0] << 120) +
      (dst120[1] << 120) +
      (dst121[0] << 121) +
      (dst122[0] << 122) +
      (dst122[1] << 122) +
      (dst123[0] << 123) +
      (dst123[1] << 123) +
      (dst124[0] << 124) +
      (dst124[1] << 124) +
      (dst125[0] << 125) +
      (dst125[1] << 125) +
      (dst126[0] << 126) +
      (dst126[1] << 126) +
      (dst127[0] << 127) +
      (dst127[1] << 127) +
      (dst128[0] << 128) +
      (dst128[1] << 128) +
      (dst129[0] << 129) +
      (dst129[1] << 129) +
      (dst130[0] << 130) +
      (dst130[1] << 130) +
      (dst131[0] << 131) +
      (dst131[1] << 131) +
      (dst132[0] << 132) +
      (dst132[1] << 132) +
      (dst133[0] << 133) +
      (dst133[1] << 133) +
      (dst134[0] << 134);
   compressor main_cmp(src000, src001, src002, src003, src004, src005, src006, src007, src008, src009, src010, src011, src012, src013, src014, src015, src016, src017, src018, src019, src020, src021, src022, src023, src024, src025, src026, src027, src028, src029, src030, src031, src032, src033, src034, src035, src036, src037, src038, src039, src040, src041, src042, src043, src044, src045, src046, src047, src048, src049, src050, src051, src052, src053, src054, src055, src056, src057, src058, src059, src060, src061, src062, src063, src064, src065, src066, src067, src068, src069, src070, src071, src072, src073, src074, src075, src076, src077, src078, src079, src080, src081, src082, src083, src084, src085, src086, src087, src088, src089, src090, src091, src092, src093, src094, src095, src096, src097, src098, src099, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, dst000, dst001, dst002, dst003, dst004, dst005, dst006, dst007, dst008, dst009, dst010, dst011, dst012, dst013, dst014, dst015, dst016, dst017, dst018, dst019, dst020, dst021, dst022, dst023, dst024, dst025, dst026, dst027, dst028, dst029, dst030, dst031, dst032, dst033, dst034, dst035, dst036, dst037, dst038, dst039, dst040, dst041, dst042, dst043, dst044, dst045, dst046, dst047, dst048, dst049, dst050, dst051, dst052, dst053, dst054, dst055, dst056, dst057, dst058, dst059, dst060, dst061, dst062, dst063, dst064, dst065, dst066, dst067, dst068, dst069, dst070, dst071, dst072, dst073, dst074, dst075, dst076, dst077, dst078, dst079, dst080, dst081, dst082, dst083, dst084, dst085, dst086, dst087, dst088, dst089, dst090, dst091, dst092, dst093, dst094, dst095, dst096, dst097, dst098, dst099, dst100, dst101, dst102, dst103, dst104, dst105, dst106, dst107, dst108, dst109, dst110, dst111, dst112, dst113, dst114, dst115, dst116, dst117, dst118, dst119, dst120, dst121, dst122, dst123, dst124, dst125, dst126, dst127, dst128, dst129, dst130, dst131, dst132, dst133, dst134);
   assign test = srcsum == dstsum;
   initial begin
      $monitor("src: 0x%x, dst: 0x%x, test: %b", srcsum, dstsum, test);
   end
   initial begin
      src000 <= 128'h0;
      src001 <= 128'h0;
      src002 <= 128'h0;
      src003 <= 128'h0;
      src004 <= 128'h0;
      src005 <= 128'h0;
      src006 <= 128'h0;
      src007 <= 128'h0;
      src008 <= 128'h0;
      src009 <= 128'h0;
      src010 <= 128'h0;
      src011 <= 128'h0;
      src012 <= 128'h0;
      src013 <= 128'h0;
      src014 <= 128'h0;
      src015 <= 128'h0;
      src016 <= 128'h0;
      src017 <= 128'h0;
      src018 <= 128'h0;
      src019 <= 128'h0;
      src020 <= 128'h0;
      src021 <= 128'h0;
      src022 <= 128'h0;
      src023 <= 128'h0;
      src024 <= 128'h0;
      src025 <= 128'h0;
      src026 <= 128'h0;
      src027 <= 128'h0;
      src028 <= 128'h0;
      src029 <= 128'h0;
      src030 <= 128'h0;
      src031 <= 128'h0;
      src032 <= 128'h0;
      src033 <= 128'h0;
      src034 <= 128'h0;
      src035 <= 128'h0;
      src036 <= 128'h0;
      src037 <= 128'h0;
      src038 <= 128'h0;
      src039 <= 128'h0;
      src040 <= 128'h0;
      src041 <= 128'h0;
      src042 <= 128'h0;
      src043 <= 128'h0;
      src044 <= 128'h0;
      src045 <= 128'h0;
      src046 <= 128'h0;
      src047 <= 128'h0;
      src048 <= 128'h0;
      src049 <= 128'h0;
      src050 <= 128'h0;
      src051 <= 128'h0;
      src052 <= 128'h0;
      src053 <= 128'h0;
      src054 <= 128'h0;
      src055 <= 128'h0;
      src056 <= 128'h0;
      src057 <= 128'h0;
      src058 <= 128'h0;
      src059 <= 128'h0;
      src060 <= 128'h0;
      src061 <= 128'h0;
      src062 <= 128'h0;
      src063 <= 128'h0;
      src064 <= 128'h0;
      src065 <= 128'h0;
      src066 <= 128'h0;
      src067 <= 128'h0;
      src068 <= 128'h0;
      src069 <= 128'h0;
      src070 <= 128'h0;
      src071 <= 128'h0;
      src072 <= 128'h0;
      src073 <= 128'h0;
      src074 <= 128'h0;
      src075 <= 128'h0;
      src076 <= 128'h0;
      src077 <= 128'h0;
      src078 <= 128'h0;
      src079 <= 128'h0;
      src080 <= 128'h0;
      src081 <= 128'h0;
      src082 <= 128'h0;
      src083 <= 128'h0;
      src084 <= 128'h0;
      src085 <= 128'h0;
      src086 <= 128'h0;
      src087 <= 128'h0;
      src088 <= 128'h0;
      src089 <= 128'h0;
      src090 <= 128'h0;
      src091 <= 128'h0;
      src092 <= 128'h0;
      src093 <= 128'h0;
      src094 <= 128'h0;
      src095 <= 128'h0;
      src096 <= 128'h0;
      src097 <= 128'h0;
      src098 <= 128'h0;
      src099 <= 128'h0;
      src100 <= 128'h0;
      src101 <= 128'h0;
      src102 <= 128'h0;
      src103 <= 128'h0;
      src104 <= 128'h0;
      src105 <= 128'h0;
      src106 <= 128'h0;
      src107 <= 128'h0;
      src108 <= 128'h0;
      src109 <= 128'h0;
      src110 <= 128'h0;
      src111 <= 128'h0;
      src112 <= 128'h0;
      src113 <= 128'h0;
      src114 <= 128'h0;
      src115 <= 128'h0;
      src116 <= 128'h0;
      src117 <= 128'h0;
      src118 <= 128'h0;
      src119 <= 128'h0;
      src120 <= 128'h0;
      src121 <= 128'h0;
      src122 <= 128'h0;
      src123 <= 128'h0;
      src124 <= 128'h0;
      src125 <= 128'h0;
      src126 <= 128'h0;
      src127 <= 128'h0;
      #1
      src000 <= 128'hffffffffffffffffffffffffffffffff;
      src001 <= 128'hffffffffffffffffffffffffffffffff;
      src002 <= 128'hffffffffffffffffffffffffffffffff;
      src003 <= 128'hffffffffffffffffffffffffffffffff;
      src004 <= 128'hffffffffffffffffffffffffffffffff;
      src005 <= 128'hffffffffffffffffffffffffffffffff;
      src006 <= 128'hffffffffffffffffffffffffffffffff;
      src007 <= 128'hffffffffffffffffffffffffffffffff;
      src008 <= 128'hffffffffffffffffffffffffffffffff;
      src009 <= 128'hffffffffffffffffffffffffffffffff;
      src010 <= 128'hffffffffffffffffffffffffffffffff;
      src011 <= 128'hffffffffffffffffffffffffffffffff;
      src012 <= 128'hffffffffffffffffffffffffffffffff;
      src013 <= 128'hffffffffffffffffffffffffffffffff;
      src014 <= 128'hffffffffffffffffffffffffffffffff;
      src015 <= 128'hffffffffffffffffffffffffffffffff;
      src016 <= 128'hffffffffffffffffffffffffffffffff;
      src017 <= 128'hffffffffffffffffffffffffffffffff;
      src018 <= 128'hffffffffffffffffffffffffffffffff;
      src019 <= 128'hffffffffffffffffffffffffffffffff;
      src020 <= 128'hffffffffffffffffffffffffffffffff;
      src021 <= 128'hffffffffffffffffffffffffffffffff;
      src022 <= 128'hffffffffffffffffffffffffffffffff;
      src023 <= 128'hffffffffffffffffffffffffffffffff;
      src024 <= 128'hffffffffffffffffffffffffffffffff;
      src025 <= 128'hffffffffffffffffffffffffffffffff;
      src026 <= 128'hffffffffffffffffffffffffffffffff;
      src027 <= 128'hffffffffffffffffffffffffffffffff;
      src028 <= 128'hffffffffffffffffffffffffffffffff;
      src029 <= 128'hffffffffffffffffffffffffffffffff;
      src030 <= 128'hffffffffffffffffffffffffffffffff;
      src031 <= 128'hffffffffffffffffffffffffffffffff;
      src032 <= 128'hffffffffffffffffffffffffffffffff;
      src033 <= 128'hffffffffffffffffffffffffffffffff;
      src034 <= 128'hffffffffffffffffffffffffffffffff;
      src035 <= 128'hffffffffffffffffffffffffffffffff;
      src036 <= 128'hffffffffffffffffffffffffffffffff;
      src037 <= 128'hffffffffffffffffffffffffffffffff;
      src038 <= 128'hffffffffffffffffffffffffffffffff;
      src039 <= 128'hffffffffffffffffffffffffffffffff;
      src040 <= 128'hffffffffffffffffffffffffffffffff;
      src041 <= 128'hffffffffffffffffffffffffffffffff;
      src042 <= 128'hffffffffffffffffffffffffffffffff;
      src043 <= 128'hffffffffffffffffffffffffffffffff;
      src044 <= 128'hffffffffffffffffffffffffffffffff;
      src045 <= 128'hffffffffffffffffffffffffffffffff;
      src046 <= 128'hffffffffffffffffffffffffffffffff;
      src047 <= 128'hffffffffffffffffffffffffffffffff;
      src048 <= 128'hffffffffffffffffffffffffffffffff;
      src049 <= 128'hffffffffffffffffffffffffffffffff;
      src050 <= 128'hffffffffffffffffffffffffffffffff;
      src051 <= 128'hffffffffffffffffffffffffffffffff;
      src052 <= 128'hffffffffffffffffffffffffffffffff;
      src053 <= 128'hffffffffffffffffffffffffffffffff;
      src054 <= 128'hffffffffffffffffffffffffffffffff;
      src055 <= 128'hffffffffffffffffffffffffffffffff;
      src056 <= 128'hffffffffffffffffffffffffffffffff;
      src057 <= 128'hffffffffffffffffffffffffffffffff;
      src058 <= 128'hffffffffffffffffffffffffffffffff;
      src059 <= 128'hffffffffffffffffffffffffffffffff;
      src060 <= 128'hffffffffffffffffffffffffffffffff;
      src061 <= 128'hffffffffffffffffffffffffffffffff;
      src062 <= 128'hffffffffffffffffffffffffffffffff;
      src063 <= 128'hffffffffffffffffffffffffffffffff;
      src064 <= 128'hffffffffffffffffffffffffffffffff;
      src065 <= 128'hffffffffffffffffffffffffffffffff;
      src066 <= 128'hffffffffffffffffffffffffffffffff;
      src067 <= 128'hffffffffffffffffffffffffffffffff;
      src068 <= 128'hffffffffffffffffffffffffffffffff;
      src069 <= 128'hffffffffffffffffffffffffffffffff;
      src070 <= 128'hffffffffffffffffffffffffffffffff;
      src071 <= 128'hffffffffffffffffffffffffffffffff;
      src072 <= 128'hffffffffffffffffffffffffffffffff;
      src073 <= 128'hffffffffffffffffffffffffffffffff;
      src074 <= 128'hffffffffffffffffffffffffffffffff;
      src075 <= 128'hffffffffffffffffffffffffffffffff;
      src076 <= 128'hffffffffffffffffffffffffffffffff;
      src077 <= 128'hffffffffffffffffffffffffffffffff;
      src078 <= 128'hffffffffffffffffffffffffffffffff;
      src079 <= 128'hffffffffffffffffffffffffffffffff;
      src080 <= 128'hffffffffffffffffffffffffffffffff;
      src081 <= 128'hffffffffffffffffffffffffffffffff;
      src082 <= 128'hffffffffffffffffffffffffffffffff;
      src083 <= 128'hffffffffffffffffffffffffffffffff;
      src084 <= 128'hffffffffffffffffffffffffffffffff;
      src085 <= 128'hffffffffffffffffffffffffffffffff;
      src086 <= 128'hffffffffffffffffffffffffffffffff;
      src087 <= 128'hffffffffffffffffffffffffffffffff;
      src088 <= 128'hffffffffffffffffffffffffffffffff;
      src089 <= 128'hffffffffffffffffffffffffffffffff;
      src090 <= 128'hffffffffffffffffffffffffffffffff;
      src091 <= 128'hffffffffffffffffffffffffffffffff;
      src092 <= 128'hffffffffffffffffffffffffffffffff;
      src093 <= 128'hffffffffffffffffffffffffffffffff;
      src094 <= 128'hffffffffffffffffffffffffffffffff;
      src095 <= 128'hffffffffffffffffffffffffffffffff;
      src096 <= 128'hffffffffffffffffffffffffffffffff;
      src097 <= 128'hffffffffffffffffffffffffffffffff;
      src098 <= 128'hffffffffffffffffffffffffffffffff;
      src099 <= 128'hffffffffffffffffffffffffffffffff;
      src100 <= 128'hffffffffffffffffffffffffffffffff;
      src101 <= 128'hffffffffffffffffffffffffffffffff;
      src102 <= 128'hffffffffffffffffffffffffffffffff;
      src103 <= 128'hffffffffffffffffffffffffffffffff;
      src104 <= 128'hffffffffffffffffffffffffffffffff;
      src105 <= 128'hffffffffffffffffffffffffffffffff;
      src106 <= 128'hffffffffffffffffffffffffffffffff;
      src107 <= 128'hffffffffffffffffffffffffffffffff;
      src108 <= 128'hffffffffffffffffffffffffffffffff;
      src109 <= 128'hffffffffffffffffffffffffffffffff;
      src110 <= 128'hffffffffffffffffffffffffffffffff;
      src111 <= 128'hffffffffffffffffffffffffffffffff;
      src112 <= 128'hffffffffffffffffffffffffffffffff;
      src113 <= 128'hffffffffffffffffffffffffffffffff;
      src114 <= 128'hffffffffffffffffffffffffffffffff;
      src115 <= 128'hffffffffffffffffffffffffffffffff;
      src116 <= 128'hffffffffffffffffffffffffffffffff;
      src117 <= 128'hffffffffffffffffffffffffffffffff;
      src118 <= 128'hffffffffffffffffffffffffffffffff;
      src119 <= 128'hffffffffffffffffffffffffffffffff;
      src120 <= 128'hffffffffffffffffffffffffffffffff;
      src121 <= 128'hffffffffffffffffffffffffffffffff;
      src122 <= 128'hffffffffffffffffffffffffffffffff;
      src123 <= 128'hffffffffffffffffffffffffffffffff;
      src124 <= 128'hffffffffffffffffffffffffffffffff;
      src125 <= 128'hffffffffffffffffffffffffffffffff;
      src126 <= 128'hffffffffffffffffffffffffffffffff;
      src127 <= 128'hffffffffffffffffffffffffffffffff;
      #1
      src000 <= 128'he3e70682c2094cac629f6fbed82c07cd;
      src001 <= 128'h82e2e662f728b4fa42485e3a0a5d2f34;
      src002 <= 128'hd4713d60c8a70639eb1167b367a9c378;
      src003 <= 128'h23a7711a8133287637ebdcd9e87a1613;
      src004 <= 128'he6f4590b9a164106cf6a659eb4862b21;
      src005 <= 128'h85776e9add84f39e71545a137a1d5006;
      src006 <= 128'hd71037d1b83e90ec17e0aa3c03983ca8;
      src007 <= 128'hf7b0b7d2cda8056c3d15eef738c1962e;
      src008 <= 128'h1759edc372ae22448b0163c1cd9d2b7d;
      src009 <= 128'h8c25166a1ff39849b4e1357d4a84eb03;
      src010 <= 128'h966e12778c1745a79a6a5f92cca74147;
      src011 <= 128'hcc45782198a6416d1775336d71eacd05;
      src012 <= 128'h4a5308cc3dfabc08935ddd725129fb7c;
      src013 <= 128'h79fdef7c42930b33a81ad477fb3675b8;
      src014 <= 128'hd7ab792809e469e6ec62b2c82648ee38;
      src015 <= 128'h467437419466e4726b5f5241f323ca74;
      src016 <= 128'h5b7c709acb175a5afb82860deabca8d0;
      src017 <= 128'h30bcab0ed857010255d44936a1515607;
      src018 <= 128'h2ba4b180cb69ca385f3f563838701a14;
      src019 <= 128'h38018b47b29a8b06daf66c5f2577bffa;
      src020 <= 128'h12f175ffae3b16ec9a27d85888c132ad;
      src021 <= 128'h176ea1b164264cd51ea45cd69371a71f;
      src022 <= 128'hf87f43fdf606254131d0b6640589f877;
      src023 <= 128'hade9b2b4efdd35f80fa34266ccfdba9b;
      src024 <= 128'h2e2950656fa231e959acdd984d125e7f;
      src025 <= 128'h98b33c6e0a14b90a7795e98680ee526e;
      src026 <= 128'h3308fb2e642aad48fcfcfa81b306d700;
      src027 <= 128'hc470f0e7f76fbfb83412fc12ac322c12;
      src028 <= 128'hd86dbf1128805c5dad1b8f60c9e4dab2;
      src029 <= 128'h2cc0f859aa6524ab713b7e05ebe21368;
      src030 <= 128'ha859890cd670f668637e0edc5b6e4ae7;
      src031 <= 128'h32f06cab0d9c2aa8f837ef727460f22;
      src032 <= 128'hbd30291a55fea08e143e2e04bdd7d19b;
      src033 <= 128'h9c31d9b25a2b745b7b59051bf40048d7;
      src034 <= 128'h983631890063e42f14aa451ca69cfb85;
      src035 <= 128'h3d4a5d5128fafd04559b5975b2d650af;
      src036 <= 128'h6a1689addfe1b30791725f0aac7c8803;
      src037 <= 128'h9145de05b3ab1b2cdf26f51766faf989;
      src038 <= 128'hbf9c0efb5816b74a985ab61c5adf681;
      src039 <= 128'hb3969057425cb200105ada6b720299e3;
      src040 <= 128'hfa83ada4a2121ac5f689a4a5ffda0336;
      src041 <= 128'hfca055362169df82b9bdee2dd663049d;
      src042 <= 128'h6ae04d52adb328cbf3158c0c66dd7794;
      src043 <= 128'h4d6b234fdfa7c6ed32d1f81ba636425c;
      src044 <= 128'h19a5711b2ea60b99fa7ff8bfb044284a;
      src045 <= 128'ha0acf4c9658de17eec3aa314da9bb017;
      src046 <= 128'h41a93f90dc8215271da3b7e2cad6e514;
      src047 <= 128'h27896389df3277fd1d77ce4058d87776;
      src048 <= 128'ha68e88e0ad4041504c14982d9ead926;
      src049 <= 128'h6f790959a3e04b3b756b0715e7180322;
      src050 <= 128'h353545792da44da189b5b368df14c612;
      src051 <= 128'h2371ea2c0247145f4a814d53964ddb77;
      src052 <= 128'hca24be4d56672017555a40854578bab3;
      src053 <= 128'h29f2c3c74505f4f60a8c46c709215f4f;
      src054 <= 128'h5c6460364a1eb1b7955d0e77fb5eb866;
      src055 <= 128'h4b1cb8bd2130260c8c69778ffd42f697;
      src056 <= 128'hef0a81ed3d5d60bcbb0378eb7a62722e;
      src057 <= 128'hd5e73e3f673617d94d7bd307122411e6;
      src058 <= 128'h57f98d1ecff4c56bf9ea2c64cc417e7c;
      src059 <= 128'h7f6b8793b318ad4c1db2b4527aa56a18;
      src060 <= 128'hceca2ee310da8a9516408169a38d8afc;
      src061 <= 128'hfa7ee0538974df5bff773ce32b2c492;
      src062 <= 128'h379deda1ade6c5e9b6e355f695bb440d;
      src063 <= 128'h2aa50f4ec6f0093395d1805142cb6d1d;
      src064 <= 128'had4ab155c09fcd8f739cd488869bdbd2;
      src065 <= 128'h41a8a6e165e049937f411fed1e70e799;
      src066 <= 128'h1ac902ee25777cf09f9821883744da64;
      src067 <= 128'h856f3d95e0ae1a1b6c596216ae0fdbc8;
      src068 <= 128'hd17034ce51797350e6256403bf3df0bb;
      src069 <= 128'hdfde228125fb5f3d866d7002091472ad;
      src070 <= 128'hd7a3283c27e969e2c8bf23fb9a431f7a;
      src071 <= 128'h10fc9eee0a1727f7ea5f24b6de6fec4b;
      src072 <= 128'hdca5b35354a1d50572d6bc20d80d6a1c;
      src073 <= 128'ha7f5195cde62d43f261908b9ccf719ab;
      src074 <= 128'h92e94e89089b30a0809f292387a1798f;
      src075 <= 128'hbf391fbb138c3460fd938adc99a2ecb1;
      src076 <= 128'hf8e45086ca819c6fd872298c7b72590b;
      src077 <= 128'he2a01335a83023ab053e4b42cc4da021;
      src078 <= 128'h6238d0a0cf5e9ea362584ab368777bab;
      src079 <= 128'h209818d1ef7e85eca417956f29ee7f3d;
      src080 <= 128'h5582a3bdd476fe38babd4745497e9f1a;
      src081 <= 128'h6af944e07b38785b0932f5b6f11ddff7;
      src082 <= 128'hc0a59677579501a62fda854775e0ec3;
      src083 <= 128'h52daad326c00984c734bb05788c31f6;
      src084 <= 128'ha145789921f8c1569e0df45b992a34a1;
      src085 <= 128'ha6245b598c94af98b3386c3e1af4787f;
      src086 <= 128'h306aa871feef71cbc915d113dc45488d;
      src087 <= 128'he6ac9d8a4160ff927c7550f20a3c2c6f;
      src088 <= 128'h254bf7ae1d0ab994f20b575d4e28e674;
      src089 <= 128'hec41e6f66c0be55c90e639e1e44fc3a9;
      src090 <= 128'h101bb5fa6a6776231ad1daaaef8d9ff0;
      src091 <= 128'h40a978bfb8f8903b53125ffdf655860b;
      src092 <= 128'h2d8b5b41590e83da586f1721078548d7;
      src093 <= 128'hd1aa6c5e3b019fcbf96d4403d48c93f3;
      src094 <= 128'h24aeba79e4b8298798ba0f0e120d7126;
      src095 <= 128'hbf7b68ae1f8941b6e6a1a40bf031f4b9;
      src096 <= 128'h2452bc39dbf2eed13b9cea959ad7558f;
      src097 <= 128'he5ce0ca6606821d6280a07ee4ec985ff;
      src098 <= 128'h390a9016cdec85da200f7753f217faac;
      src099 <= 128'hc13e66af3c9590d33e2aad3e82221345;
      src100 <= 128'ha9c72e7b6b770df15f59aa2c4a82e06a;
      src101 <= 128'h542bd7599e8c82821da132cdc68d4fd;
      src102 <= 128'h21cc14b312bdf75fb3c161c313f2a37c;
      src103 <= 128'h877a2133f2ed33e1a31559405e87905a;
      src104 <= 128'h70f8dd9952177eb7e6b920daba6a098f;
      src105 <= 128'h788c161ef3cc9d8a4b1678e45f20f406;
      src106 <= 128'h1bce35d8cbe88a3f2f7a304ff344c911;
      src107 <= 128'hb02de52c9b050db28ee4fd021cb66f67;
      src108 <= 128'heda2fc4c7237d420b3dd77e1cbb02fe9;
      src109 <= 128'h6e84f8ea6bf4d047c4841a8d2f751bde;
      src110 <= 128'hc149fa8e7bb8c2f11624d318a32652e8;
      src111 <= 128'hb2f11ef9d48644820078cb124b7350d1;
      src112 <= 128'h37fef6b501fda698764657ca9e65736c;
      src113 <= 128'ha100ed14fa92cd28c4c536fb1d4d1180;
      src114 <= 128'had9d1f4217b18e6e78aff58ec058a332;
      src115 <= 128'hfbe86a8ea1cf0d1d47b3df4167c21355;
      src116 <= 128'hab2212c9e23b580e4523dbbb1eeed219;
      src117 <= 128'h71d04b0f656fa7e6b5c03f6f94e4cc44;
      src118 <= 128'hcad00273120961ea0913508715d38ca9;
      src119 <= 128'hdc66a27b6a325333116e8a6429deb984;
      src120 <= 128'h1af55c2688083ebc35d4cd35a08c3a00;
      src121 <= 128'h47534952c9c5fef1e76f8a76c74f11cd;
      src122 <= 128'ha0f9c0749177b6d45f2e9167713eceb1;
      src123 <= 128'h1eda4209b270af551f9078d52835bcdb;
      src124 <= 128'ha1d20ebc5aa3892a4c88b9d8ab12fb53;
      src125 <= 128'h7a0a02ba37cf80256a447a90be0a5a56;
      src126 <= 128'h4cd8ef2471a8c9c60f6ab75bf55b2e5c;
      src127 <= 128'h78b61daf5afb9565068a3c383739076a;
      #1
      src000 <= 128'hddfae808afd8643211035083fa999f9b;
      src001 <= 128'ha8aa1e45c7cbc6201a4f7a165264961;
      src002 <= 128'h92a651d7c069c542240397213a082921;
      src003 <= 128'h54a8762b2b12c92c62565a955487b5c3;
      src004 <= 128'h6f6ddf79affe2554e5aef699a5e3a719;
      src005 <= 128'he90f79f835783f662114c2d650ea1324;
      src006 <= 128'hfbc59e92ca1209ad596305b371b221e4;
      src007 <= 128'ha217cf253be957670884fd16636abf8c;
      src008 <= 128'h7552c6e86953a1155a62ddc4e2091f49;
      src009 <= 128'h7460d20d94b9cdb56e3c18c9ef1fa0a3;
      src010 <= 128'h3725bd0c79c45c38b440ffe0413770e2;
      src011 <= 128'hd7422560b36f3cd0acfeba4441030ae;
      src012 <= 128'ha795ac544a30f7cd00fdec23598ca3b4;
      src013 <= 128'h315e80807425f4e93891aef5ebe0572c;
      src014 <= 128'he2014a459b3a0c891a32e1489bbac838;
      src015 <= 128'h8930d17952ab793f51abf5e5cb775e24;
      src016 <= 128'h14827a895e6364c630ac79dd0b5aafef;
      src017 <= 128'hdc2897c6845398134fee71444d236555;
      src018 <= 128'hcf1accc1eaca38110c26e5d9702dc88a;
      src019 <= 128'h70aaf52575e417dd7e5b637dfa98c115;
      src020 <= 128'h2e2dffdff57b8a920a12f3b364fc0dba;
      src021 <= 128'he64ddd918e9b185e1b770deb6f51ea78;
      src022 <= 128'h42d01ba3a2652c9e89421c6d764ab510;
      src023 <= 128'hbb9e5a022c2df3c219518f87b63f83c6;
      src024 <= 128'hcbdc014dbedb42e6da313e783e9973b;
      src025 <= 128'ha91da2cd8bf06f64b4178592b76fc5b2;
      src026 <= 128'he6cd3595d4f0d65dbd6817b638b80611;
      src027 <= 128'hacb5959f4eb9876884a5b1c31095e497;
      src028 <= 128'h7af2f402a0e624f15f89d54d3bcd6aec;
      src029 <= 128'hcf4bb31523254d812bdfb7279501e917;
      src030 <= 128'hc3d9b3b022b56be11392a255fdc12930;
      src031 <= 128'h36a52df9f8247e70b2194ff3c46ac0d6;
      src032 <= 128'h974d9d499bc698825a7c831a62759469;
      src033 <= 128'heaf94919e69b79717f9b76efa1057256;
      src034 <= 128'h4f06ea1874a264447d3c279b5bce228b;
      src035 <= 128'ha71b80ef8e36b82f3856be31f568c9c6;
      src036 <= 128'hd25ab04930e9be17b413420866dfeb1e;
      src037 <= 128'hf19b43da6253dfe34aaeb212c90ded29;
      src038 <= 128'hdceb201357d9af8d3fe65f90f631681e;
      src039 <= 128'ha867a0f0a8e6a772b9cde60cab1e6794;
      src040 <= 128'h298e9a79abecfc0b581ba30742965873;
      src041 <= 128'h8a1d8b4292d6ff735b3a4595045892c1;
      src042 <= 128'h5a79b46a26b61b06a1645f58bb78eb2d;
      src043 <= 128'h649def50fb2de1ea0b976c27db931ce;
      src044 <= 128'hff9d318d22a3a621109197853a081a6;
      src045 <= 128'h6f6a219672ef7dce376e22a6ec071cf1;
      src046 <= 128'ha629d3322d4ba5a44fdc13515ba830dc;
      src047 <= 128'hbf4fa4a3c90853fdfc9ea692ba626aee;
      src048 <= 128'he413961f68c6dd5e027752fe61f68c6e;
      src049 <= 128'hc253763876703835b476998dafc8128a;
      src050 <= 128'h8024532000cbd3132bdb572063eaa07f;
      src051 <= 128'h1463c5f825ee54abb3191702bb80d98d;
      src052 <= 128'hd216ad53d4088ff7d71330613cc4f772;
      src053 <= 128'hb7c144fb2b16ad048fb87c76af044a8d;
      src054 <= 128'h990e8f01dd5aacc7ed7a6edf6d5b7d50;
      src055 <= 128'hb5c99b49751f7e54a0e774869ed9c124;
      src056 <= 128'h40a210150a40a3799a1ab3579d6c84af;
      src057 <= 128'h606375b8bb937826bcee9d29ce4f1ca0;
      src058 <= 128'h94c0230e3b4df81eeb3462ca032149d;
      src059 <= 128'habf0f4bd4af0a6fe5bbdd1f416f14aad;
      src060 <= 128'h5b1654ad81e774de3c740119754724dd;
      src061 <= 128'h566ff3ec679b29e8c0c32da9bc49b58e;
      src062 <= 128'h6480fdc0f1c58f447e083c1bcda6a326;
      src063 <= 128'hb8acdd816522ff4674b7061c09ce15a8;
      src064 <= 128'hd18533e7efa2faf58ba0bf3675e0c52;
      src065 <= 128'h8c626a9fee4e6bcbd6deb9245e695b1;
      src066 <= 128'h8429aeae877e5ea1c33993f235045f77;
      src067 <= 128'hf8cc3f3bd59b148ffa7bff5f62d59938;
      src068 <= 128'hfb52451d90e7e1a11db1dfdc357f0a64;
      src069 <= 128'hecadbb86f16f1487f7f21e5cce0755e3;
      src070 <= 128'hd0fce92295be263b0253dc8cd1f0c570;
      src071 <= 128'h583678eef3ca5f6427fa8b8a909b471c;
      src072 <= 128'h52b049944b1dd9fda02ebb764a8b77da;
      src073 <= 128'h300a21879cb9f9aabf4ddeaa41f2005b;
      src074 <= 128'h2b7bde99878f40ed2c805ac7d48457df;
      src075 <= 128'h94665d45284b7bcda3af11d0a8ab29f1;
      src076 <= 128'h6f446806c1378e75627b9de79ae445e0;
      src077 <= 128'h8df7a26786fadb0e89b1e0d44218ca25;
      src078 <= 128'hd840fccb2446eceecaa0a6796e83a7b2;
      src079 <= 128'h903374bfc81236e6ec77cfc8b38e5adb;
      src080 <= 128'he65a3ae43a72017dc29ed120cddb2316;
      src081 <= 128'hf0fcccc6fb46ed398772c3475cba9be3;
      src082 <= 128'h3df8eeefe44a01f69251ad083fcb34fa;
      src083 <= 128'hed2ee36fc2112edaf1e7ea9b2f6570d7;
      src084 <= 128'hec6e61bd70c455a92a1bc11230331476;
      src085 <= 128'h53e836639c14940d5b2d81ccc602bd20;
      src086 <= 128'h65dcac6cc329870a33e9e55e402492a3;
      src087 <= 128'hd2928f4be1514a0db27516ea63a6aae9;
      src088 <= 128'h4741ee56b5e2834d907d85322076d932;
      src089 <= 128'h12677895c6be59658f16c91dd6d47e4;
      src090 <= 128'h67fece7f1ff06dcf45aa79bd855fb35;
      src091 <= 128'h29b496640f52361d82f1240d4e5c6dd2;
      src092 <= 128'hb93c2989c399fd7fb75db71ea4531fe9;
      src093 <= 128'hb56b9357b34dc8b053f3c15842ce91c0;
      src094 <= 128'hef7dee1a8476af98425de95fc846bf90;
      src095 <= 128'h83210210a43c991d2d4da4ef95e38180;
      src096 <= 128'hca8033a7a5fd89c831610b3d1257363c;
      src097 <= 128'h8e50c79ac582644479faf5012287401b;
      src098 <= 128'h848610cfd21276c21519401c8b1f1137;
      src099 <= 128'h147a08acc65d8e4ed01e488b00a1402e;
      src100 <= 128'h91fd7d4a5a31a6a69b87cc5e6d7fe9b2;
      src101 <= 128'h832c9b7960c8e5a0d560e64c55f7792a;
      src102 <= 128'ha2f62516dc88b09cd7604342fcbc3229;
      src103 <= 128'h5d156b6eceec38d511fcda922d80170;
      src104 <= 128'hcbf8e26a4fae667bb2e74e770fe1cedf;
      src105 <= 128'hdd35d11688181a813d1ea49ed469bf4;
      src106 <= 128'h2e4025346987b05274219d3ecdc39412;
      src107 <= 128'h18a775945b8c4949106861d3633d9c54;
      src108 <= 128'h2d5590c90576598359cd012a06b42b6f;
      src109 <= 128'he5a1bdaea747795eb0c952af9db31510;
      src110 <= 128'h79fe0a1b7efbe877b1e186d7df254e5d;
      src111 <= 128'hdcb32e4a891dfa7b0d3dc6aadba45b5e;
      src112 <= 128'heceb9505dbc33e56c8a17945ca6d3e06;
      src113 <= 128'h8771fe6f7d870b678ac870419365f61;
      src114 <= 128'hce03a34da022dfee843fb606e8b7e2da;
      src115 <= 128'h606e8502002f9cc4096bfafff5b7751f;
      src116 <= 128'hb22b89748c5c192ff1c51dda28280370;
      src117 <= 128'hebbe1a41c781e11f2cb38568291a58af;
      src118 <= 128'hf212cc6f540988e79fed6060ef23d4af;
      src119 <= 128'hf75a7e6f2b863694541d1a814815642c;
      src120 <= 128'he0db22d329e316ad39ddc4775a220eb2;
      src121 <= 128'h90bccb66e06314505d0057167680891b;
      src122 <= 128'h3729e33c5507d2b909e7f7862f25291;
      src123 <= 128'hafdb4e0b01716f1d956a2f20ee283bb7;
      src124 <= 128'hfff83cec2c05b870cd34bcd7b7ed75b4;
      src125 <= 128'h18b7f1a2f74f190559c07423a89f5916;
      src126 <= 128'h789c3c723ee29e686fa00319e54ce0de;
      src127 <= 128'h94d50a99eba0842465a5ac1f7b2ecfc5;
      #1
      src000 <= 128'he072caae797c27bfc79385209c921e7f;
      src001 <= 128'ha0483bb2f6d080c46409df32cc4e66da;
      src002 <= 128'hc78c2f9da418b24e0acf9ff88d3281a;
      src003 <= 128'hc48ae37406dc1579647640a1b6a659ef;
      src004 <= 128'h64a2bc48f9fb4010dec772b7bb22fa31;
      src005 <= 128'h572abb532b6b7b42295023267644d183;
      src006 <= 128'h80e97f74c30759a448a133abdd55daaf;
      src007 <= 128'h956c2129b934718f2d492ca241f4317d;
      src008 <= 128'ha9d499ca2698c2d614f1ddc4bc972ce;
      src009 <= 128'haea6231508ef444a6e63ffa48d2ad974;
      src010 <= 128'h354af1bdba5612f7600aa45e44e1b08c;
      src011 <= 128'h9cf600ec1c3c8d3521d4fb7e22587c89;
      src012 <= 128'h93a25c9b6e3a52d707fe6a4e2a6f1e47;
      src013 <= 128'h2b52dab12367ad9e8dcd7d64b9e8e4ee;
      src014 <= 128'hd68d2bc2dac7c336ea045534f6796fd3;
      src015 <= 128'he63317c3430342c7dcfbde0ac5fee487;
      src016 <= 128'hf7f1bb2780665563a0c30ce957ac59f2;
      src017 <= 128'he983cc1d25033a3eb1f5d7d0887b4cca;
      src018 <= 128'h8e33dcabbe684e2bbd637b3afc0b1519;
      src019 <= 128'hfe1c51e5ea31e67ae16802053c0a94de;
      src020 <= 128'hfef06b0468fc642af6f259264e60678b;
      src021 <= 128'hf924e06aaef5baef1903b45fd01cf935;
      src022 <= 128'he47516941d8ac1a902af33820938ad77;
      src023 <= 128'h517fa07e7b0f78c1b8f35c26d13ec39c;
      src024 <= 128'h2b02237ee2cd159aebba80d2820bc51d;
      src025 <= 128'haf04ef81b5481bf2702cebbe3544f189;
      src026 <= 128'h67ba6b1a96954911a4e0ee5b1638325c;
      src027 <= 128'h749d4601df98377981bd53363bac2660;
      src028 <= 128'ha51de78b8d00b7b27d82fccf81eb88e5;
      src029 <= 128'h74f8c57b24c582caeab3c4d8d4e4004b;
      src030 <= 128'h179d221d8e5f37fa68f49b51f3fa8613;
      src031 <= 128'h1c622f82d0813d923aca43f27b777bf2;
      src032 <= 128'h181a218ecfd645605c05c1f3241d3e27;
      src033 <= 128'h32d116fe8f08963c962488052305e6d3;
      src034 <= 128'h8f3e64f479140a61ee65afeb1b674518;
      src035 <= 128'hdf61c53457d1d37cc7afae8fdfecb2ae;
      src036 <= 128'h3a05c0b73ddf55b2015128dbaf8c96a9;
      src037 <= 128'h4642cddb4fbe2aaefbf70946d6ada066;
      src038 <= 128'h17776c3a57435d9ced3032ed824c6948;
      src039 <= 128'hef96a21449b3fe663b4c0730253df737;
      src040 <= 128'h1e94eb4bc74f73cad4c667bb211e55c3;
      src041 <= 128'h78916712de5fe0ee801095005ae52530;
      src042 <= 128'h277dfc7b722c353d1ee1723b4a9686a4;
      src043 <= 128'h3a8be1617fd2770a568d6f3ef4b445aa;
      src044 <= 128'h6382f3b5f9adf8c56247b40dae5ceb3d;
      src045 <= 128'h9e3b3f04d418864590de6fbaffb59512;
      src046 <= 128'h4fab2ad88091a21d6637c09facf606fc;
      src047 <= 128'haf157ed9849648e85084a40f3b8f5fc7;
      src048 <= 128'hf7b37a86d21dbc093a357442f325f875;
      src049 <= 128'hc57842a9934c472a0c72fe13fbf28c1c;
      src050 <= 128'h88da091b61f6c8770212585b0b2f8580;
      src051 <= 128'h6a4ace0ed89a95009f13d2fbe583847f;
      src052 <= 128'h3bfb255eed0d04182d58bce989745cd7;
      src053 <= 128'hf45c88409da283380a8bc856c3edd9b7;
      src054 <= 128'hb42fb35758d97f4a95331356074f3be0;
      src055 <= 128'h1790a6b7845c21e7988d0e4a2266a107;
      src056 <= 128'h1a7e256db6ffe12c1a6f0c9af1f7e90f;
      src057 <= 128'h339fbb6951cd2c07a8f78b61f9d2b2de;
      src058 <= 128'h8f41d3e41eceb5e5801841f4820d15c6;
      src059 <= 128'h2dbdb6e57844c2ac729bd820e4ad24e2;
      src060 <= 128'h6a8d3e8420fe652b56fe23018c3af69e;
      src061 <= 128'h816480fa90a2b8e1141bd89660924d2b;
      src062 <= 128'h3bcab3eadcff697dd26d028dd1f15ee7;
      src063 <= 128'h6df2fc823956fba972323dc9c67781b2;
      src064 <= 128'h241813ef799fde337a2be04940d2d16f;
      src065 <= 128'ha73e3f3b5c27761d4894d9fc70df67b9;
      src066 <= 128'h166a1a98af3b5a9185bab545d4e26a5b;
      src067 <= 128'h27b51ee70f1a6c44f239fbb01f6ceec1;
      src068 <= 128'h77f63854e668bb6ec408143f290d07e4;
      src069 <= 128'h7f00625769560c063008a519ad830951;
      src070 <= 128'h855a7d8dd46e34aaae9d1797c284e0be;
      src071 <= 128'h86c976870fe3cfc991ab513369fe284;
      src072 <= 128'hd7f14ec29a9dadd2e7aad0707cddb4cc;
      src073 <= 128'h21b6323246b7d9bb2966398e4a295d;
      src074 <= 128'h5690f74daedab7b5e2aa55a7495103ed;
      src075 <= 128'h702a5b67b7ae77585b45cf5ad7de701d;
      src076 <= 128'h258694b6113c183677f4531bfde9d47d;
      src077 <= 128'h3513198c67f8ab5705727bb50bee2ebd;
      src078 <= 128'hab341860fefd320bf5efaa99010f5ddf;
      src079 <= 128'h7d5d9031e80bb7eba49999cf87e51bbc;
      src080 <= 128'h10e857f88986148f8b3e00e76151787e;
      src081 <= 128'hbeb9c9e2156e3ae54fe4b7355c29b6da;
      src082 <= 128'h773b83502743e0df5e15428a833cf90f;
      src083 <= 128'h61f9c40838330558fb2323e7d6a2c379;
      src084 <= 128'h56fb5c72ed6a1bfc81be81f4bef874d7;
      src085 <= 128'hef82c4d6438dc8b1971964f8d2fb05ca;
      src086 <= 128'h51c6a2e46f48744f7abc9f0b86fe0ded;
      src087 <= 128'h1dd95d4c0637fdcadf4630adbaaa6300;
      src088 <= 128'hf64e8f4aef89c2e7aa1706669b6e83a9;
      src089 <= 128'h7f79ee0e299cb482449213ac2fab184;
      src090 <= 128'h1d8cca3b6261479043a061c445a16970;
      src091 <= 128'h8d5f52c083f0ba7756b8002a0f424ffa;
      src092 <= 128'hd1cae1937ed61f4ee875176629530a13;
      src093 <= 128'h54e27ea64202faf9dcebef56a31ca36b;
      src094 <= 128'h961139cfffbdfd47dc7972f0133894b3;
      src095 <= 128'h662701363aeb5bc0f63d307ca9d21bf8;
      src096 <= 128'h706146ffbecba4c8b2c92c129bd91220;
      src097 <= 128'hd4062cce773a13fb37503d7733672754;
      src098 <= 128'h8fce7af52c1b3c7f33c4233c833b07e;
      src099 <= 128'hcda840fd4adb0798039d60ba9c993735;
      src100 <= 128'hfaa2cbad467a6bdfb63c1dd82a9e9a38;
      src101 <= 128'hdd7516f558aa03838dff06d28340fed5;
      src102 <= 128'h2c94151d52fa3935ff28355076847398;
      src103 <= 128'hd5e32aef05dd1ef0080638c9496749fb;
      src104 <= 128'h49954cf1faaf500ca74b3d208c3fa29f;
      src105 <= 128'h6b291a13637c3644c9345ce70e5bc44c;
      src106 <= 128'hf367dbe240e3469f39b66d71951a0518;
      src107 <= 128'h6c749cf41f7550bcb550f22172e55360;
      src108 <= 128'h7d5e121623a35ae7a31a27cced4dd7c;
      src109 <= 128'hd3100ac51932263c4eec95b014c30b50;
      src110 <= 128'h700b1433f5d6147620f12d46e775f27e;
      src111 <= 128'h86861f295cb76bb9c0ff34b4e4bd7d57;
      src112 <= 128'h7ff5101d3f1cd31b86ff76d11fe32b56;
      src113 <= 128'h5b7801ea86343347daa6b26ae30d04fd;
      src114 <= 128'hcc869dea38a7ac5426b1caba3fccb2c1;
      src115 <= 128'h2e665ecb06f9f4e68b4eb003401a2e8a;
      src116 <= 128'h2826ef27f190cb53b489f5c7e22f6e82;
      src117 <= 128'hbeb778d62b021118ae63ad3a94d7f681;
      src118 <= 128'h697b85380ff73f2533251c76d8efb5c9;
      src119 <= 128'h3665b6a5634da412816a5ea8618a4763;
      src120 <= 128'h1a608f0d7e4132ad86b0915a8880f9fd;
      src121 <= 128'hbee5f64d3e37355efbdc678abf33551d;
      src122 <= 128'hfc145cfe469a1289ac91c01e734c5192;
      src123 <= 128'h65739938a96e2bf4586523b8f9154865;
      src124 <= 128'hc315d334e47c98ea139e5ca2b9e7f780;
      src125 <= 128'h723dc8f5b17078ee112930f2cf21ae6a;
      src126 <= 128'h992e7dea037432634a0609aa827acd0d;
      src127 <= 128'hdafd518dd55f0e0eef6be029bbef627f;
      #1
      src000 <= 128'h793910e656e16c2b659badcb9bcae27d;
      src001 <= 128'hd197b56179b68b9523aa9e6770bc3ec1;
      src002 <= 128'he9bf79f4b3739067cf085288f0041e32;
      src003 <= 128'h9a642c24a34acc3eda68fa2a59581c94;
      src004 <= 128'h3055d84e3c38bfd6d7e239089090d244;
      src005 <= 128'h4d3903626ef4d6b4424c222f577aa515;
      src006 <= 128'h41ca37f5f7de1a6131bf3b36bac114b5;
      src007 <= 128'hdfa2e52bd35169bc0044c690f17a7c84;
      src008 <= 128'h9e3f4f152f5c5cbee55b88fff0862962;
      src009 <= 128'hdec22e0cd4cd82fa2adfd824edaeec39;
      src010 <= 128'hdbb59fc25cffc96ebd03c81f7ff35029;
      src011 <= 128'hc8359b916e935faf9502e1d5167ad089;
      src012 <= 128'h2c14af79c4a0c1cd0654f465b311d9c4;
      src013 <= 128'h624aadaeebbcf1f6dedff24b3567c813;
      src014 <= 128'h2dc6c2accbae0e932f39c04551bb91c1;
      src015 <= 128'hb425aae7eb533c3a0879fbdc7843b3;
      src016 <= 128'hfa2225d77c6d8ae1463e4336bf3cfe56;
      src017 <= 128'h832e9e1e1b908d6de5e6190b28da2b89;
      src018 <= 128'h9ba66e98679140e0b6fece9a8f15c995;
      src019 <= 128'hc99d5f9ec634effdf02dd043d01acef6;
      src020 <= 128'hd6b6b5d01c87284dc5fa8ac995a37efe;
      src021 <= 128'hc3ac232caf405e52199a1949ba9d82b8;
      src022 <= 128'h9b9a9bf50a78491f0211550313218ef7;
      src023 <= 128'hb3f175d015c7a82023f3e5aed1de4fa8;
      src024 <= 128'hfc7aad95bfdf8a9e9446d493a4d6ce54;
      src025 <= 128'h8bdd4b9dfc2cd5c7d5562dabf4a9b4e3;
      src026 <= 128'he6e4ac85f10185fd8f81598725394778;
      src027 <= 128'hf49eb5a696ab64d235128906a4ed017b;
      src028 <= 128'h7837e5069398dbd616db36e4d4ae3486;
      src029 <= 128'hdcbcd86ea2e86f7add6af484024d65de;
      src030 <= 128'h81de9808c2ff347bd527b331240eb6c1;
      src031 <= 128'hf4098aef1d50fccffec09878f0344058;
      src032 <= 128'hc045883b940f737e548c3ec425365ca8;
      src033 <= 128'h40fd8aaa3504e26c5f7e07d3160d0b9e;
      src034 <= 128'h50c6735014b3f2641598734a86c52c1b;
      src035 <= 128'h8ace37d3673ef518c6cbb1796239f30a;
      src036 <= 128'h8d17e6327e8aeae24a703e3120a202f;
      src037 <= 128'haa0cc3271daa42fc90b15e3da5005582;
      src038 <= 128'h4d7e444990b6e394448236e9863c6992;
      src039 <= 128'hba13834fde8e3228aa648f16f0355088;
      src040 <= 128'h808ea422c6f6d1d53b77ba5f586076e3;
      src041 <= 128'hfa29559dc81a58a66245b749b9a6edc1;
      src042 <= 128'h1c3df9183278f64cae1367a579e9b08;
      src043 <= 128'h1c67556d79acd84313b2cc1593098549;
      src044 <= 128'h44ee50715745ef5a2e0885fc5da23c06;
      src045 <= 128'hb9c3a78fc8d3aceed370c51fd8e2ba4c;
      src046 <= 128'hbd2098c6c2de59500b2f72efec0959b8;
      src047 <= 128'heda04e30ff741d1ca8936bd386a29efb;
      src048 <= 128'habbebd4ff9e590e4d36d8076998b1e1c;
      src049 <= 128'h9411723a50b417eb7111f1d19c8fe812;
      src050 <= 128'h832cb6a724e2e13aa0e5bd8cdd7524bc;
      src051 <= 128'h61880ea05e5ecd0a3cbafcaa643580a0;
      src052 <= 128'hf66b72a94142452b361c57ab3d992624;
      src053 <= 128'h257ea412a21574899fbd4b9f56756682;
      src054 <= 128'hc2862234d81580dc24d878a13e5aed83;
      src055 <= 128'hec023a99e4c80a291d5f9dfc98b0b4d7;
      src056 <= 128'he79d1be27f29e86c8a730eaa16bb4fb0;
      src057 <= 128'h8301c5b945ffa36b63c2523d4b32bc86;
      src058 <= 128'hf4e35152312cd4340b177efd054f0566;
      src059 <= 128'h806094aa4037fffa14b8317e75555ded;
      src060 <= 128'hd05d2cb96b76911f7c8765b6b04a2620;
      src061 <= 128'hf08502ee47e3d101d72e0feea289858;
      src062 <= 128'hea8760aada4dda766a34bfb4e62a3fb5;
      src063 <= 128'had283c0df230400a386b01c05ffe6c11;
      src064 <= 128'hfd6cc3648191cbeb175bf448a0ce5b5f;
      src065 <= 128'h835875c3952049e4a8fcf210dac15a07;
      src066 <= 128'h3c241ca590425d14e6b0643c188417d8;
      src067 <= 128'h39dc2c06f38075439722bf902f073516;
      src068 <= 128'h42045f8c3a72a669e03cc361214e10ee;
      src069 <= 128'h96bad500ded1b80232e977612e975c72;
      src070 <= 128'hbdc5a588d0ab9ea4c15f47ca204e6817;
      src071 <= 128'h208d549b6b0efd0100dd28b3acea35a3;
      src072 <= 128'h80d9a24e0a83303889de7a2c7c26c722;
      src073 <= 128'h2ca5f0cbab78a4ee385127f1f317930e;
      src074 <= 128'h714d85bde1976c14aa069b5b510d115a;
      src075 <= 128'hbbe74e1ba3289b58a62f45c2f0cc8eec;
      src076 <= 128'h19b2b59530519f6ab51e3a7bacdf3038;
      src077 <= 128'h60252b8d2cd9f51a10c313bd6478a399;
      src078 <= 128'ha6d5eb2ee891f80c970a06dcf444adae;
      src079 <= 128'h24e9031675f80092ea4f44cfeafd080b;
      src080 <= 128'h89419b16bbca76e0e56a47e742f81126;
      src081 <= 128'hbd335a642d79f3f6ca92720ac2e8fae2;
      src082 <= 128'h53b9a632f967522170c4340643db0235;
      src083 <= 128'h8e7a744a7f3c30f26e5e2da91b92f8b;
      src084 <= 128'h77fd7fd135cb60f26a75e179fd14f9d4;
      src085 <= 128'hac69c00681b84ea71f21747566f0f769;
      src086 <= 128'h8439ba12afd65c3a7484ffbbfd9de84;
      src087 <= 128'h9937f592185aeb983d9f3e803ba68577;
      src088 <= 128'h37ef373e32dec6d586901942366e3cca;
      src089 <= 128'hdbf9a793ecb9cb393103d90417426bd0;
      src090 <= 128'h9efb00b7a397b217851143e593aae480;
      src091 <= 128'h7647513c9e6e6309a553472a15b74ad;
      src092 <= 128'hc9d4e1bbc4d3fec2faf3d90e586a7302;
      src093 <= 128'hf9873b5e08dfc975a4fd9204b3b9e84e;
      src094 <= 128'hae9e8d0384983111371a239070c742d0;
      src095 <= 128'h3c91e45824b27e8301cbd9c2d35f581e;
      src096 <= 128'he1289e96ebe3387b68cbaa9e22d72fab;
      src097 <= 128'h486cf4d67c23bbfc0490642fdb5bf01f;
      src098 <= 128'h82042c0b1da221b825454e29ad5ac10c;
      src099 <= 128'h135981c7b984dbe3aef82d2e51f83e44;
      src100 <= 128'h310dfbf4d7418ae8cfa71765e757155d;
      src101 <= 128'hb2835bff857d114b4b91cbe8fea4ca6a;
      src102 <= 128'h60fc01e2bcd635ccb9c4abb6a6a99aab;
      src103 <= 128'h13bd01ae70dd4704248988cf091523be;
      src104 <= 128'h86d6c42427b22a70a9452a96a1239c72;
      src105 <= 128'h599490667d4165889a347cdad4814f7f;
      src106 <= 128'h92976e6ce04d350f260aeef295dd24bd;
      src107 <= 128'h2997e8996059c8a9cb0206728fff6a1a;
      src108 <= 128'h848d77e3c7975813ba4e199cf2b8fd15;
      src109 <= 128'hdf302d42c4545268acc08d9899dfd2f5;
      src110 <= 128'h478947081b08fdc11162ce262d64584a;
      src111 <= 128'hfdf0d6056b7b2370940ca324420a746a;
      src112 <= 128'h5536212a58d776da0f013f4e73961f8e;
      src113 <= 128'he7d37bcc63f6ed2d68652c4da322e658;
      src114 <= 128'h3deaf9a0a724dc8f4be669fbfbdc2233;
      src115 <= 128'hb888cb6597b19d4f16d24a67c6b1b41f;
      src116 <= 128'h368712c085dc1819df6316b93f739143;
      src117 <= 128'hfcfd32468884b81da7e1572891c9992f;
      src118 <= 128'h184dc5184c596a49334f97a4ec8bd978;
      src119 <= 128'hc66456bfe73ce3cc4306dd16a5b466b4;
      src120 <= 128'h732f3e8b251bf7645e302bed15ade79c;
      src121 <= 128'h72824622a4b0c73bf74e21a162e5b726;
      src122 <= 128'h847eabd3be5c193391a69f34d7cbd7ff;
      src123 <= 128'h444c3c0601ed02dbd6638406290af021;
      src124 <= 128'h41d1240bb53c902262885f8cd6fb2221;
      src125 <= 128'h7f562e989bd23ec521f943546776eb37;
      src126 <= 128'hb1a8e5c62c075d2cdf9e407af3531a52;
      src127 <= 128'ha85536f31bf8fbebd06e62e6dc5a2a83;
      #1
      src000 <= 128'ha416c71df64d977c20a4ef0eee68e406;
      src001 <= 128'h6fb5545cd95cd1ae6d7cefa55aa2356b;
      src002 <= 128'hfc8847d21b067b10958620855d587077;
      src003 <= 128'h218a6b1873ecaee9cd00f4288ec14f83;
      src004 <= 128'h7ae1a24ea792b2b462e1b434b3670f54;
      src005 <= 128'h18bcaa21b887d3e9a317105664afbf49;
      src006 <= 128'h86def5a0474fc1f74d26c0c52ba08a24;
      src007 <= 128'h565e5ae7ad82e067ab3594148ed2b26b;
      src008 <= 128'h17d9fa660063b5c924fa9196f8015987;
      src009 <= 128'hd8cd5da373cc35245675f2fcc0ca3f4d;
      src010 <= 128'h1a6ed97f03cd7bab667b94c973213530;
      src011 <= 128'h352d6f27b98713be5462a18d1b6d6ce9;
      src012 <= 128'hc736e1668042e02f1d7322518b763f63;
      src013 <= 128'h2a1fff41af1b70131c7bc6c8d62fee8c;
      src014 <= 128'h8f8b36e406fa11b492294b0bd4ed425f;
      src015 <= 128'h19b6b91b1f695a01f5f5b0d2042e4fec;
      src016 <= 128'h61a5c06ec4be5a7fa15d41c915369965;
      src017 <= 128'h3ac2496e62436476b9298df641a97327;
      src018 <= 128'h5f1fc0aa486998f52d51d8b76579644;
      src019 <= 128'hd0fe4a59329ec4ac2ea5cef8e6b724ce;
      src020 <= 128'he08aec96f4159113cac4b9e6778d028c;
      src021 <= 128'h912d791d3288a67e030c98e85e2408fa;
      src022 <= 128'h9d0a4fac67aaa0688dcfb198f0e51f30;
      src023 <= 128'h9ddd6df0329b638600bc698bea264afb;
      src024 <= 128'hfb813983106fa2ec4896c62cb397b350;
      src025 <= 128'ha4b2f62c610097fb589c25911608f0df;
      src026 <= 128'h487eb3df3b71e722c579009ca3efb3de;
      src027 <= 128'hac606a5d49dd3b0ea29d06e06f5714d7;
      src028 <= 128'hd31470c8acb14314662a7671276d105c;
      src029 <= 128'h99c5e64cb8c6773e9610c047f84907a1;
      src030 <= 128'h4dd6862a5ea2fdfb8c33cf4d783d4a6d;
      src031 <= 128'h6ca992350989e9e258beb6672b8059d7;
      src032 <= 128'h3b2559fb54d6aa2dfd7fc7de3a0cc176;
      src033 <= 128'h27ef096756bf5e579ff9b0f506274afb;
      src034 <= 128'he0934e387f42af90e412eb0bd260a30d;
      src035 <= 128'hfd577ceaa623c2783a94f14b08302ee6;
      src036 <= 128'hacd85b9f6ff00a21add7ae79eb0f6c21;
      src037 <= 128'h70bef8fb659812bf4a18bafe2df4a748;
      src038 <= 128'h28ce122009b12bc988054048f53a7cec;
      src039 <= 128'hbba6ad3cd094d2af793dd40f1de16841;
      src040 <= 128'h4d433c1f4e25a42bcc4589b5bbd4b4ed;
      src041 <= 128'h44672c65d1e0a50e9602634b08453d3e;
      src042 <= 128'h4b3099ecd4364172b60b7264a69cfd32;
      src043 <= 128'ha2334974746c8933eee69c71ee166b74;
      src044 <= 128'h1cf7f935e6cc9e41768599decffd101;
      src045 <= 128'ha939e190c6f1c3ad9b86d80d10b8c060;
      src046 <= 128'hef38123719a0f532d2197d9333a70c3d;
      src047 <= 128'h1a143f918a34065b2b058a0ee3531771;
      src048 <= 128'hd9836a1fbad8ae6a5f5ce777dae3c720;
      src049 <= 128'h9ade0a942709483a176f9018b18646ce;
      src050 <= 128'h816241bd5a57cde5f13fc40b489b9a03;
      src051 <= 128'h24a3b63500513063020aca12055dfed4;
      src052 <= 128'haaa91ed47be1251abc1255417d534839;
      src053 <= 128'hd13d78bc42c07c7ef7402ba246884eed;
      src054 <= 128'h52d1de24bf3ba58ed02fe51359eea30b;
      src055 <= 128'h4056125ca1ddc5a325053d917eb78350;
      src056 <= 128'hcc9bd78e5a456f863e3292dbb0bd6bdd;
      src057 <= 128'h8eace752634ad5b9fd72a908edb8a483;
      src058 <= 128'h3b48146954fe81bba3455904083087b4;
      src059 <= 128'hfb20fab5be98e6d20bf2e1da430e055c;
      src060 <= 128'hada6b225c607fad901fe2e706aa066f7;
      src061 <= 128'hb56ac802c76f432cdc5aa6c9d1abd865;
      src062 <= 128'h2bc38de01d0820e0a24921ff8616ba88;
      src063 <= 128'h1541c1e420fedb80ae9e2e6adaa21ca;
      src064 <= 128'h54536cba289f88b49b566e06cc800b04;
      src065 <= 128'hf77b8c86ea3249e632ab7704d185cd3a;
      src066 <= 128'hf634dbae9e7be7ad97d8c97d731b8cf9;
      src067 <= 128'h5d7ee6e358bdd490d26c34f8f6b1557e;
      src068 <= 128'h6b35da2c04465ea7cabf5c57c5795b58;
      src069 <= 128'he6ab5199de9318967ada5a662fa0823a;
      src070 <= 128'h7e8c83ecbf9582c79d592226302d6194;
      src071 <= 128'h916b3d918b55fde8968a9f2884eee7;
      src072 <= 128'h2f40d4efbfb553c2fd162e6fe93cef4b;
      src073 <= 128'h2d26904840131e33277b20adfefed218;
      src074 <= 128'ha5160d17e71f767485883d4441b11180;
      src075 <= 128'h6ca1c7a8ba71d93589d9a4015207cce5;
      src076 <= 128'h9af1b4564034dca41eb6217876cf14a2;
      src077 <= 128'h48ef09a4b8c0ace840a0864341cb57da;
      src078 <= 128'h808b20f6f281e24c8384841da56a4a75;
      src079 <= 128'hf7243a0c0947bf82b8ed3aa4681be70b;
      src080 <= 128'h683e8e1cfb99a06b6649e79473b8bf6;
      src081 <= 128'h9b6f338a0665be98c138418d964ede98;
      src082 <= 128'h111244066e30d1ba4ed0081835d2cfcb;
      src083 <= 128'h9b39285ec9cf17ba2a51d1ea18eec8cc;
      src084 <= 128'hef1a030cfba98e7520f37df2a0fe1900;
      src085 <= 128'hfdeb26efcced6bffb92f5f3d86634e4a;
      src086 <= 128'h2539021523c0b46981001b5e21366a11;
      src087 <= 128'hb5560b631cef5445707f76cef137c97;
      src088 <= 128'h14b92ea4421f4828902a94ca22a85558;
      src089 <= 128'he1b9f50e216d9a63eb8313a85b53cd42;
      src090 <= 128'h547008340af23ed35ee10379e9afa682;
      src091 <= 128'had5a14c79fce833719c613bae1bd8bab;
      src092 <= 128'hdad389fe6af26631176151c236c55e3b;
      src093 <= 128'hab5c31226e9393387c7e8bd2f19348ca;
      src094 <= 128'hcf31d2c4125b65b14483cf58312bccf8;
      src095 <= 128'h3efc91f057f599d1732ae464cf762ef8;
      src096 <= 128'hb473e51420a7446bf9c8d852760eff62;
      src097 <= 128'h2783662b7f49db7a38168876cda5a0a0;
      src098 <= 128'ha9333123166533672c97f169516bb4ed;
      src099 <= 128'h1cc99fcc1ddbb059ffb9c71bb69d0fae;
      src100 <= 128'h4f47bc9453e6db96c24507885272898f;
      src101 <= 128'h6287fadd330a90c317310ddb2101c5;
      src102 <= 128'ha3b0cc064d6bbd5da64b62d5a889ea84;
      src103 <= 128'h28b671b88eca745cd90f6bbc2b7513d8;
      src104 <= 128'hb484db42e58000cf427585d8e5379893;
      src105 <= 128'h16d91fc5be85039460fc74e80d0d82f9;
      src106 <= 128'h1cf0589debde3e110ec5c62d24020912;
      src107 <= 128'hd370bdf9d85d37fe4d5866cee64f0edb;
      src108 <= 128'ha06d8653567494dfc399daf6444ef491;
      src109 <= 128'h842f9c6554fedaa0173e585cd5b2fd55;
      src110 <= 128'h4d628581ff6dc856c9e93ebecc0afa36;
      src111 <= 128'h5961640123d8c4800e67287ccf127621;
      src112 <= 128'h3b2d1fc9eded54e339e6f58f7fdf2229;
      src113 <= 128'h70a22d8ec3c02b36ea727bf4202aae64;
      src114 <= 128'h3985577fc069f48d5c5815b0197aef97;
      src115 <= 128'h4bc61ffdc61053ed451b1c8ce0c012d2;
      src116 <= 128'heab5f50a9f2a5843af3357209f7b8a2e;
      src117 <= 128'h70910cca4fd0fda21c32a1ded54f58b7;
      src118 <= 128'hdec0efbf60339ee9a8b12ccabcc0cdcf;
      src119 <= 128'h567ffb07cbc968749bb3aa4c5147a3fa;
      src120 <= 128'h7e8fed3dfde60dd454b3f5c1ff9e16ef;
      src121 <= 128'hd83dd24bbcd8d4e4b8d056c18506b30c;
      src122 <= 128'hce5e761b7b59a1c0bd08b032f9ad5202;
      src123 <= 128'hd98efec68fdeab3c158423a5005ba4e1;
      src124 <= 128'hdf0644a8c3d7df292368db81da34effa;
      src125 <= 128'hacdb9ccc100dcfdbc413b8e8319c7b43;
      src126 <= 128'h6b3190f4e55ef7495e3fafbffc06d3de;
      src127 <= 128'he2cd813001e1dd8c91a7859b39147d0e;
      #1
      src000 <= 128'ha2d9281b94334bb0103ba901337faf64;
      src001 <= 128'hc9aadaa6e440aa7ce95361bfee628c9a;
      src002 <= 128'h860e7019579dc1fb73d0c8bfe2fb8f04;
      src003 <= 128'hc176eadbe5173c41fdf156226751d1a4;
      src004 <= 128'hc0b2ae8b77887200b6bd58d6e8c2215d;
      src005 <= 128'haeb405f1d006434cedb52ad7db3d977b;
      src006 <= 128'h7a31daf12dcbb10ef7a15f3beb5dc17d;
      src007 <= 128'h81992dc5d7488a7680aaf97e454b57c1;
      src008 <= 128'ha94f30d62f595bc0dad16c2b96561c94;
      src009 <= 128'h3f848dfcefd622d77b3402f41f13fea5;
      src010 <= 128'h975e2ac2f08df7c1e20fed4b182f0297;
      src011 <= 128'ha5660feb35b996bd901d169d25ab3477;
      src012 <= 128'h606d396e18867eb5199121865dbfc02b;
      src013 <= 128'h49777f5b9a614ac871a953e291f1955c;
      src014 <= 128'hfdfcbce0d6fdf5166b1a37c623ed6d79;
      src015 <= 128'hb016dddaecb501ee2d8cf7e121583621;
      src016 <= 128'h531d07a1ad26ebe4cadf4be2468f6365;
      src017 <= 128'h657475fd1720b8b4c12c9c8d199c4745;
      src018 <= 128'hed1a474854b58fb5cd656a213f8beccd;
      src019 <= 128'h10c565d554059bed1fb861a396d53ecf;
      src020 <= 128'h3eb913924c041d5a7e41b9af9ba78849;
      src021 <= 128'h584957f20f1f41f3b6ec93b4df0b60b9;
      src022 <= 128'h8f72b28c16fca750fa679a042b44d7a2;
      src023 <= 128'hdb3d663628e1a8afa02255129ed03a7e;
      src024 <= 128'h913e7095fff706948ecc8c9dbc0f91ee;
      src025 <= 128'h4881f40077dd23074593b102f9ae8048;
      src026 <= 128'h71d6ec10cceeba877d3c106227d20e84;
      src027 <= 128'h27bcb21ae8497caa531bbb0e9be82d6c;
      src028 <= 128'hd9f415ff4c786b1e06d341c5ceb885eb;
      src029 <= 128'hcfc76634cea323b493df0c5af3afc368;
      src030 <= 128'h56eebfe7f5a182c5d246fd226b8f76fa;
      src031 <= 128'h151a3787d03e6d922b243c589743dbc8;
      src032 <= 128'hd8821713e97a194e6ef93741721e4596;
      src033 <= 128'hbeb6533abca281f1c1c7f10be0467889;
      src034 <= 128'hcd024ec04b2bac3c5950d2bd900e7701;
      src035 <= 128'h47f559efb76db463b9f15b792d53f13c;
      src036 <= 128'h1e682c1ff26b659bf85cfc9ecf130e07;
      src037 <= 128'h6966437363eca19aed3696ce2f914af5;
      src038 <= 128'hbe0d894c52f29d2c3747414b1140e8ae;
      src039 <= 128'hf95b88a89600a0436bbde06429a8f86;
      src040 <= 128'h267ce9c1166fca8f91627297fdf3aece;
      src041 <= 128'hca6838d1cec5aed28b9d2bd6d88cf5ba;
      src042 <= 128'hcabfcd948beace4de4f440284f4f2f74;
      src043 <= 128'h92ecd51d031e3c424dc557e294ad6516;
      src044 <= 128'hf685b1f354271488122594275aa27950;
      src045 <= 128'hd219c7785891a706c43b5096d39e4b11;
      src046 <= 128'h5a23c2f2262acd409067f7264ce68c93;
      src047 <= 128'h22b62906685b54ed17d4cc0e8bb1f29;
      src048 <= 128'h91fd78156e3f32e8d22428c03bc3f21f;
      src049 <= 128'ha77e6a1dda6d27207a1cfb21b85e81d;
      src050 <= 128'hd4055fa2d660600a0c35a424a158972b;
      src051 <= 128'h3335219c09224fa0365d3eed327bb556;
      src052 <= 128'h631c3308c3007cb168f76fd638d34dd6;
      src053 <= 128'heb4194a05cd65445d05366ccb051460d;
      src054 <= 128'h3a4bcaab8659cf439de8ddf4a4b10a7d;
      src055 <= 128'h1c6d0e358a5082e214079f9eba95b4f6;
      src056 <= 128'h73665614da72eb92a4be525e134e7a5;
      src057 <= 128'hca1871c69e7b6789873c6d8bfeeb9881;
      src058 <= 128'haa88496556547b4d317588ff44296fe7;
      src059 <= 128'h7df8b7f044a1d4d0d6dffc21b1c2ed56;
      src060 <= 128'hfee2f56b0ee1ce2b4b385492d4c6700b;
      src061 <= 128'h48e003be5bf2b6a11b95cd28b2764173;
      src062 <= 128'haf5f7bd63021c8ad3302a5cad4ae04b3;
      src063 <= 128'haf56d7ba6f086f6588df03070b320459;
      src064 <= 128'h2c8941bd4b7118acc2411753bd3a98bd;
      src065 <= 128'hccfcd7467a440b3413e34b3d3d946990;
      src066 <= 128'hee51bca044c0a5ed6d2db46a5bb955f9;
      src067 <= 128'hc490758166ab247a75fe000cc40732b4;
      src068 <= 128'h4fc3489b9c14c815d24f8f4351a2fa15;
      src069 <= 128'h97ec1a4076ad98ba10fb5581cccb4dfb;
      src070 <= 128'hde6ff3f11ce76bc0c34c3f471171c294;
      src071 <= 128'h1b742111a032943c4ab878c73b342529;
      src072 <= 128'he8d7025b8a8bc03efafd02b84b990ee7;
      src073 <= 128'h3f74df9ae43bd5309b3e660550835669;
      src074 <= 128'haeef4b09bc7838b31a9af2a3ec6b2ea2;
      src075 <= 128'hb5ed09cc8320446942493187676b94a1;
      src076 <= 128'he771edcc969a2550fdb9def338428c7a;
      src077 <= 128'hd4323934cda9cfae10ff4de8e6ff73b5;
      src078 <= 128'habe04a6109ca574d20979829cc898b6a;
      src079 <= 128'h7194a9f14114fa1055b3b1acc34920a7;
      src080 <= 128'ha35c56b352403e1dbb8bb9ae57e061c6;
      src081 <= 128'hb7d52dcef2aaaaf0e8ebbae25bc1c77a;
      src082 <= 128'h6f1f7a150631d91b5073039f1e6ad906;
      src083 <= 128'hf6bd16ac4ab507018e6b81a3e9edc59c;
      src084 <= 128'h10a15299054efa504962073ba0f9986a;
      src085 <= 128'h61af473df106892ba1fa46f346685cdd;
      src086 <= 128'h73f19747e9a28f3cb9abe19f2911cf30;
      src087 <= 128'hcb771b1e922ba0aae055b94fdcb8a6e;
      src088 <= 128'haaf5cc090de68b59c48418135eabd8f7;
      src089 <= 128'h415fd4f37f137c0d39e65a53dd59195f;
      src090 <= 128'hc68ddf7dd7d5f9bdd3e47e37817d6729;
      src091 <= 128'h1b04eaa423f33d55192489473b6b8130;
      src092 <= 128'h6f0667649d672b49cdbdc97fb9fddad9;
      src093 <= 128'hf9646b27b465260092c47c9950625b3b;
      src094 <= 128'h446781798383818fb235872ff68273bd;
      src095 <= 128'hbe3bcc6457446b2dddb3d8ee6f8b6cbe;
      src096 <= 128'h96bead62d52da285543e882cb7068b26;
      src097 <= 128'h4aec0bdee2f75b1efda59820148a3cf;
      src098 <= 128'h439c6004ebfc2aa5c8c7e9554d27653e;
      src099 <= 128'h9a7945cf66c10396be8809a6f1e902dd;
      src100 <= 128'h54bb58bd4e8b1b517a0cd3b5e85c7c1b;
      src101 <= 128'h4b5e5471c640070899d80fa6f0f4c87c;
      src102 <= 128'h27503d1e1756e0d4b187594d577b1f95;
      src103 <= 128'h5942adbad0576ddf43237e0874d43d6d;
      src104 <= 128'h4251bdb2776adad8744f957ff7d9dde9;
      src105 <= 128'hc68b1f6e0d5e1bd98d8320312c2747c0;
      src106 <= 128'h551a9eb6dcade3bff755b4635c340e94;
      src107 <= 128'h5759b929ab9873c46246ce0a0e9920ec;
      src108 <= 128'h79e32aa0e2238f5548e422fdf89ed0ff;
      src109 <= 128'ha0766bc39ecbcf97c201af5a45276f0f;
      src110 <= 128'h9d930454e6219ba45be01ab72c7db93f;
      src111 <= 128'h77c6f07dba43cf43b1aaafb1d1958c;
      src112 <= 128'hf77bf1ce58fb42053e7498a7286334df;
      src113 <= 128'hc33cedaa40c0ab3dfc753aa1d0f64d2;
      src114 <= 128'h530d9dac09650fe0d5df6c49994269b4;
      src115 <= 128'hf7a2b187758eff25033f692fad9d81e7;
      src116 <= 128'h77183b112d130744b253a6353652e007;
      src117 <= 128'h231e58b01acd382443ab4db80e45aea5;
      src118 <= 128'h95999d257b4b57fe556133371177fc2c;
      src119 <= 128'h61f35552d1576498ada375ee049167c9;
      src120 <= 128'he0db4322f8b8b8b5863a5de90aea39ec;
      src121 <= 128'h8fb91db81d3b7cfbbd317f2fb72d9bb4;
      src122 <= 128'hb720fabacc5d5cd8265244e8501de827;
      src123 <= 128'h7e6f85818a6993de7e10b8849271c546;
      src124 <= 128'h2c05fec343305aa1725b40ca2e001a75;
      src125 <= 128'ha05206d25774a8f0bc7300c9d918cda4;
      src126 <= 128'hf26093e5ae1c4447c43097a8e212335f;
      src127 <= 128'h993c47c3f953249aff29867d22c0f031;
      #1
      src000 <= 128'h4f567492a3ee0dd9054a516e5007181;
      src001 <= 128'h23b982e5141ba7b127a917799450826f;
      src002 <= 128'h6391a567684e8ede2fca7a048c39ceab;
      src003 <= 128'hc50613abc67518c95e19d2bd028f1175;
      src004 <= 128'h109122085d81778a5ef70581af71f4ae;
      src005 <= 128'hec85a655c8a8135a816db439d2a679ac;
      src006 <= 128'h2a5debfa9dd0630e189798129ee3efdb;
      src007 <= 128'h7257d90043240b2d77cc7a7b4162ca27;
      src008 <= 128'h18ef618f5c4250886b28d7d6651bf718;
      src009 <= 128'hca82007fdb0b921f426afb9c2653b39e;
      src010 <= 128'h14b64d4fc5483917729730a1560e409d;
      src011 <= 128'h95099cd0285f9f8a33213ea434f956f1;
      src012 <= 128'hc3ee79d13e85bc2ab4095a99962cd344;
      src013 <= 128'h70eb1aee07e53dfc22f062975d96425e;
      src014 <= 128'hfef89ac90d5e0895d7511fe6183fc86a;
      src015 <= 128'h3306f416b09b81639ff67b314a15d941;
      src016 <= 128'h9d02e44cb5e5f25ddefa351400c99f27;
      src017 <= 128'hfa0ab3567b113deedeeefbd673ce1e6;
      src018 <= 128'hd493227edcd3c1302ad735da2d11b499;
      src019 <= 128'h7303ca039f7642908104908f1f32140f;
      src020 <= 128'h5048b85ac544b042c9e6358375273ef4;
      src021 <= 128'hc17fe224820df53f591eb142dd4f1ac3;
      src022 <= 128'h75029fbd561d047914d277e4ff0f84c;
      src023 <= 128'h34fef75045709961232d7ed8b2192894;
      src024 <= 128'h9f95ecca4972e2d0dcdef04303f9c3a3;
      src025 <= 128'he90a23643a03873ebb9bdf46f5930c38;
      src026 <= 128'h9bef38facbce125bda1c0162387e3cae;
      src027 <= 128'h8dc118edcd492f0c93c6023fa2b24fd9;
      src028 <= 128'hfce10181e6bac20520168140c55752ec;
      src029 <= 128'hd3f1e7dfa84cd94a656f075e99691df6;
      src030 <= 128'h247b34f7cc2c158b4f46089758500c02;
      src031 <= 128'hf25dcd20ee526cf5ced15cd37641cd98;
      src032 <= 128'h86d2660533d69c6168f8a67abdf76a13;
      src033 <= 128'h1a8f1af06ce2ecf9dd295d4db0b03350;
      src034 <= 128'hc10b89c02692a85929bfce744531ff00;
      src035 <= 128'h58dbc60f29f123022160af294ead1428;
      src036 <= 128'hcc9546b397cd20ac93b21689df84f6fb;
      src037 <= 128'h489782b2495f350593247ace409c3af1;
      src038 <= 128'h42b42bf869e5ab7b1b9c26485f000fa2;
      src039 <= 128'he7bdcaccf1d04cc8eb0f052f003abfe;
      src040 <= 128'h9b7f3e1b6c953dddba85eeec576b3230;
      src041 <= 128'h6cdd497d1e8be9c33a98eb14cd1fe22d;
      src042 <= 128'h2044eeef025e816b0a53381b267739f7;
      src043 <= 128'h7370a76cf8af92d5d73b293d2eaa2c7;
      src044 <= 128'h8dc73e489e293bd91ae3b6381c723c20;
      src045 <= 128'h8e106701a478856a52a068f73613b453;
      src046 <= 128'he644d4f4e0985dd30a813be624f1b0a6;
      src047 <= 128'h5abd752ea30047d0085d7943eb63d7ef;
      src048 <= 128'h56a0da9e350a2abc695d5d5a1da8f429;
      src049 <= 128'h85b535edf5d6f87902eb8a14340ace11;
      src050 <= 128'h8263da78405087bdff555ae5553da58a;
      src051 <= 128'h90eee95136487b1e944846ec7fb032ec;
      src052 <= 128'h1bb19aa0a9392defe7cc081690f089f3;
      src053 <= 128'hc82dd85819f8b828a40aaab86ea4e398;
      src054 <= 128'h190be786fe27a780f7b2b3d74873d80b;
      src055 <= 128'h7aed04c4643d87ba18c2a569109d5b97;
      src056 <= 128'h21653fa639989ec0531d32b6e80c5c54;
      src057 <= 128'h91fdbb38b6e2d1e40a22b2ce234e85fe;
      src058 <= 128'h8d40d5428c0f53727a03ee5c77b9611e;
      src059 <= 128'h736243ad72fd518f1a1d81de4b9cfdfa;
      src060 <= 128'h431c327f6e15039a59cbdf86676b9e5d;
      src061 <= 128'h3633cb67e33666a1fadc0b74f81721d5;
      src062 <= 128'h509dbfdf944e13df4a12d0df3988ba0f;
      src063 <= 128'ha4cbda9954e4960c73fa5ecd4cfec3f6;
      src064 <= 128'h1b2d8cd061c96b448e4924b8e6802d85;
      src065 <= 128'ha9fc795dc3d0db4bac9c74e2cdeb0960;
      src066 <= 128'hdf116459befa60afb0a095849ed8bfa8;
      src067 <= 128'ha161960086983739a1550300e07d5b15;
      src068 <= 128'h8a68c17bc11e95c392a55f24d592d2ca;
      src069 <= 128'h2e40d5cc1bb9967b19c87c0747951f79;
      src070 <= 128'h3d3617798dfd001027ce5dbadce4708a;
      src071 <= 128'he9f1c34d9ad02d70eb0b5d4a7baaa17c;
      src072 <= 128'hdf29a50e133d9e6fd9d7b48a7cefa36f;
      src073 <= 128'h27ca44921e51f22aff893bcfc3e3187b;
      src074 <= 128'h6b9cfa617da9c122ac2f5716df539ccb;
      src075 <= 128'h8ca5773131243f80cfedf6319bcaa8e0;
      src076 <= 128'haa07c6e1b284b450fec264ee8d6ba9fc;
      src077 <= 128'he077fb540c588f77238b0af3cf0d39bb;
      src078 <= 128'haa8c4f547ad4f768953f2ad962e5d7a7;
      src079 <= 128'h6bbd4a43cd8df058be046bc798ad2354;
      src080 <= 128'h8870582ade8204b8a3d56b4dc5c22c02;
      src081 <= 128'hd7d9cd2c352abdc0d492a3f9d7413bcd;
      src082 <= 128'h1a00cb0031f1f4f44c9dc9a84da3ea8f;
      src083 <= 128'h29f1ca3a88af77d3f15fe2ff689a0ced;
      src084 <= 128'hadfd429f70a3eddd79fb3bcdf3826505;
      src085 <= 128'h43d3c1cd44436c48cfbb5634862ac9bc;
      src086 <= 128'h6a7b14540f784eb0c966727b29af9e17;
      src087 <= 128'heca9451844587bbe0a669218613bbe30;
      src088 <= 128'h9727212f92938a3ff3c09c1aa943ccd2;
      src089 <= 128'h3c9111d08f28b6f3fc7887009dcc3e8f;
      src090 <= 128'h550a89dbb99cf8dadc016a1ee64c8980;
      src091 <= 128'ha34ac29a3f2c15697c88ad60ec35be28;
      src092 <= 128'h318f7ba99ec8c47825a65b8f44f773bc;
      src093 <= 128'hb79104d4e51e79030364180e226ed286;
      src094 <= 128'h2afebabba6f33d64c5572d91f86ad017;
      src095 <= 128'h3b6ef9a882562466b86dbb5d7650b755;
      src096 <= 128'h525bf551665c5421ec5f3b268f230a71;
      src097 <= 128'hf33131c98ec02e1bccca57a3b1eadb0;
      src098 <= 128'hcd62fd36d5f2437e95dc506c99d8adaf;
      src099 <= 128'h5dde624c6d8de017582e3ae1b812e5f;
      src100 <= 128'he777592e6f599e20400a06e95ab8a31b;
      src101 <= 128'h3ae1ab400dfe24b90d1b85c99427ad92;
      src102 <= 128'h483b995a9c834a7cb990c977f4235c2c;
      src103 <= 128'h6a33596c5684797b2a1926e5274e7c9a;
      src104 <= 128'hca4d7e3a759e9cbe6ba735b1b5f1e073;
      src105 <= 128'hbc1e8fbb61c2dec4258878d3a0a1fdd7;
      src106 <= 128'hf544412b8fb5f417de2c4c68688df8af;
      src107 <= 128'h485e5204474682516cfd088b581e00f8;
      src108 <= 128'h910f0feda2776fdff94cd0da156d3de3;
      src109 <= 128'hed6420ba3260141eb828ceb008b8427a;
      src110 <= 128'h48d44211bb047d03b1f2dfcc5dcfcf61;
      src111 <= 128'h9fe62e363162ef95096b03e621a43722;
      src112 <= 128'h4b5c31ed72bbccfc34ff496ad52583c8;
      src113 <= 128'hb94f684927ba334f90be68d55aa970d9;
      src114 <= 128'h602d808cc27efe7edff0ad7864b34997;
      src115 <= 128'hc8d13ca07dc01482c8160df50957f0c1;
      src116 <= 128'hde699e1e2922bc1d47ede52834910d03;
      src117 <= 128'h9d592a7b2542cff6071001c5c02e3a7a;
      src118 <= 128'h4c4e1314343bcd00913edb040b652dbd;
      src119 <= 128'haa757aa516daf6a65945e764b07fa381;
      src120 <= 128'h94ed072c9e781e1a394fadcd5d1ee1f3;
      src121 <= 128'ha8adc7e35bb0ecd619e3bfe6cb7033b7;
      src122 <= 128'hdf1b925e6f66be879a4c2227abac92b4;
      src123 <= 128'h84eb42d367c45071ba8a82eaad527daa;
      src124 <= 128'hfd3b748d278223ab29377d76f11ff82f;
      src125 <= 128'hdc0f71ff12ef4ae2746ddff4865d2030;
      src126 <= 128'h970ea1aac76f98aeedf3d0246f88c633;
      src127 <= 128'h119c21c47e39fd94f850cbeca7f5794c;
      #1
      src000 <= 128'h9e8be2457ad60b01efac72285dde1a4b;
      src001 <= 128'h5a0b37e8769f513a6b223250fb2d35f7;
      src002 <= 128'hb081690ac73cab38250d0c9ca556df18;
      src003 <= 128'ha7e5963c493b1112868a9123aa4b938e;
      src004 <= 128'h2e6984c6472005457b9ba35c8e296c03;
      src005 <= 128'he68f7b05e46cf2ada450d1d0d35e1fbb;
      src006 <= 128'h3fa8122d0bded21608633195e960a9f6;
      src007 <= 128'h17737931a6e49e29f7d3664bc53b6776;
      src008 <= 128'h98d0cbb77844e648601b7208f7f3032b;
      src009 <= 128'h4ae5e3ef0c5380244744ac61df73276;
      src010 <= 128'h11279e770c132eec9b1958d87961464b;
      src011 <= 128'ha31679290e618684e5a61f880c461b54;
      src012 <= 128'h7e8efd0d0279648dc8d4f7fb439e5f60;
      src013 <= 128'h8e3f4eae19b5024ceee2a362cccbcb6e;
      src014 <= 128'hfae203e1a7fd116ed8f5817f85bdca63;
      src015 <= 128'h860d23d64c85e837f5cf489783c8e374;
      src016 <= 128'h113ed69c5a8ce27b2f70b365286c6c4a;
      src017 <= 128'h1c6258f0272c763d87a60c7c41175ae3;
      src018 <= 128'hc9aaa56d0b2ce172fb4fb36eb79098c;
      src019 <= 128'h90c31d6007f1a41e8f18c17af0dd0920;
      src020 <= 128'h87bc43feff10c1d0e276b0f04551cbe;
      src021 <= 128'h53d9ba8ed3cbdcdccb650ac53bc35d42;
      src022 <= 128'h48e411b317604557b30979faf8900be8;
      src023 <= 128'hc314f367f98408a60ec003b677760e5d;
      src024 <= 128'he4ad31211c57b0c9bdfdb88eae4fd0d7;
      src025 <= 128'h5d98abc9eae9c546446c1893c9d3cdb9;
      src026 <= 128'h55e0637c7d490adf234877e301d04d0f;
      src027 <= 128'h8da28b08d71080d93bbd199b9e54afa6;
      src028 <= 128'ha04777d10efa49d4610153bdc65937de;
      src029 <= 128'h90916a5f97ad1730763cd2743719509c;
      src030 <= 128'he4e59c4ff2233a76f7bf8f347151735c;
      src031 <= 128'h9b99a16ade2523c0f987dcbc59fcd9c0;
      src032 <= 128'h1b53d85fbaaa418ba5a97fd2e2c71ba1;
      src033 <= 128'h3d3021855fbb63036c10e43363985173;
      src034 <= 128'hef6c59995f93f6e9e36b26fad9d2a060;
      src035 <= 128'h2ee6c16d351e7fc8d6ab5c68606db8e5;
      src036 <= 128'h2a05004a271fb4e55d67ed180be3fdd4;
      src037 <= 128'h527f3113f7a8992f4a058311c4791523;
      src038 <= 128'h23bae9a976c6bf55a9b932bc23500fca;
      src039 <= 128'h5a344fd7a13429cefb73ca968a5dd636;
      src040 <= 128'head6b26ab6600ef91f4e7e4c3417ccdf;
      src041 <= 128'h3affeda39c91536ba383dfb5dfc4043f;
      src042 <= 128'h3cc020d910ca65f479da713d74784fcf;
      src043 <= 128'h32a88b74992c6631e924bbb0cb8a27fb;
      src044 <= 128'hb1ddd8114c09baf401df38055f188cea;
      src045 <= 128'h69259d812a2e0ea75834aeaf0f332bab;
      src046 <= 128'ha8f7ce912532687eb173a40ae53ae519;
      src047 <= 128'h5ee97e15fedb37503714752506ce943;
      src048 <= 128'hac8d4df50eebc74086c2ae063f5bc2f1;
      src049 <= 128'h68e720101978be2860f71863ebc295a2;
      src050 <= 128'h92b8a1e10815f8138802bd32dc6b7272;
      src051 <= 128'h2d6d9fa99859792c2a865fb4eda3852f;
      src052 <= 128'h30ea170473df09482da0ca27fbda1657;
      src053 <= 128'h636f82737c16b60ae17c280b787d13e2;
      src054 <= 128'hc29e1c4f19706b9ba208bc2ba7211de8;
      src055 <= 128'he154d19d7c39c32a72916b340a648b77;
      src056 <= 128'h61dbbd3653ceaa74bc849a73f149e41e;
      src057 <= 128'h658f520cd22acfa45e9fc1a4eeb8ded2;
      src058 <= 128'h1cf922542db3c31abeca21d69570c92;
      src059 <= 128'h36feebec5df0ff7b75240e44ecfd67c2;
      src060 <= 128'haab8ef95a4b49941b231466cbb447105;
      src061 <= 128'h85505347a626ac793d8abfe328059a51;
      src062 <= 128'hfd62c146afba65cdd600b473d90d9833;
      src063 <= 128'hc61a423b2f5a140222c878274e132492;
      src064 <= 128'h4bbca2b4b54cf8e1f78441186747424e;
      src065 <= 128'h6a256d90d9e2a4c57b57619f73705a40;
      src066 <= 128'hd00b4607f5feaca1a6fee8326b63619e;
      src067 <= 128'ha0384ddf57cd8e617dcc7312db7f780e;
      src068 <= 128'hff837007113e7a58e73295ca705426b1;
      src069 <= 128'h88e985bddbebd3a4bf99cc5ed4e1efa1;
      src070 <= 128'h9fa54b2b4baf452ce107e332a64de767;
      src071 <= 128'he6437b65c63c3d085ab5d4c101a95f82;
      src072 <= 128'h816702841d62367eaf64704637ab26b4;
      src073 <= 128'h4329e4990dbf36118c9af4941e34efba;
      src074 <= 128'h969e30058225d841263d70cec5d18ed5;
      src075 <= 128'h7b6fbe5540136ca46810ae359c195380;
      src076 <= 128'h262894d153710d59b77fd039924ab4e2;
      src077 <= 128'hc2faf63731920482626a7f3ec9ce7799;
      src078 <= 128'hb6cfa3f8fc72dd60c468c13818714c59;
      src079 <= 128'h596888410df5d972076ef1af37eb9bfb;
      src080 <= 128'h4fd27dc04a4d2091733e6301f28faeb0;
      src081 <= 128'h9bd657abecb8739d87f663905f230e6d;
      src082 <= 128'hfccb11625311cb54a0665299e7f63ec0;
      src083 <= 128'h88ace67d44466000cc4c171759b5b7a3;
      src084 <= 128'hf55fdaedcf6f1f1f22fe927dae7efb14;
      src085 <= 128'hbda98d6bde047110f36418a05939ab39;
      src086 <= 128'h69223a46cdd48f958b04fdf233dc9af7;
      src087 <= 128'hfa2c00661af7ecb83e7bb18f8f13c71b;
      src088 <= 128'h7e4ab70a36e238e5a609567c4e762047;
      src089 <= 128'h5d3dc7b6fa5e8461c9e224c5780cf076;
      src090 <= 128'h79a59fb90f8320e2a3cbd5d5c05774;
      src091 <= 128'hf48a7aeb100de1140d1908c8461aac84;
      src092 <= 128'h55f7b9a0c069bfca5a3377af845c0808;
      src093 <= 128'h4dbd90c8f690304077ba5bb297d37fad;
      src094 <= 128'h5f199a64c9fd032b9d22c8861a4b1ee6;
      src095 <= 128'hc37164aa95fbda85c6c017dce8bd9438;
      src096 <= 128'hdfdade0ea9b0a8ae4f8529fcca8162d4;
      src097 <= 128'h395ad1897a40240ad297a1895710c060;
      src098 <= 128'h3796300d1ebfdb889bed02eb51a5040;
      src099 <= 128'he18a97bc913c019056b67e24ec4f4771;
      src100 <= 128'h6e3624a150fb1ee49346212ac82e7612;
      src101 <= 128'h7aefa28728dff27a30c6a6477a5d92dc;
      src102 <= 128'h60b77fae29466b49057ff1bee77bebcf;
      src103 <= 128'h750320d7acf2ad7e39b07a24c285676a;
      src104 <= 128'h866f679932faabac1c1b009e1c793cde;
      src105 <= 128'hefe23b7f412222e82e10b1a5ef9f0c0b;
      src106 <= 128'hfa35444be9aba97f8652433c94a2fc1a;
      src107 <= 128'h390cfd7e9c9da0d29087bf0e9206d547;
      src108 <= 128'h3d140b67332177e4aac8b42ceb11f63c;
      src109 <= 128'h64cb2808eae41deb9edcf3a9beb78d97;
      src110 <= 128'h2650b12408adb4a26daa3c860c2ed22d;
      src111 <= 128'h732df7ec93a27c9d050ac8ea317bf366;
      src112 <= 128'h350000267927eac4aa6fd1856fe84fa9;
      src113 <= 128'hb6c843e413250452ac29c1bfb0791b94;
      src114 <= 128'hd9249e45083a7379a850d907047e7966;
      src115 <= 128'h708e308a7875be9799fff4ba97bbd507;
      src116 <= 128'h80f2f7b17294be45deb6eee6b17672e2;
      src117 <= 128'hee95755b0a9a55983ee9ca9a4081b1e5;
      src118 <= 128'hea963dc8c05f4b53fddcfa71d52ac5a0;
      src119 <= 128'hfd04a69befb0512f3e5dcc5735397165;
      src120 <= 128'hb60bfaff9fea730f0483bea650dd55ec;
      src121 <= 128'hcd15c2fa3814553216a7276e0c9cf350;
      src122 <= 128'h8904da261b2fd815b8e32a6b990ea430;
      src123 <= 128'hcdd1e1663317f126a0cb72ad45f4eaa8;
      src124 <= 128'h2f27ae3295896e6cd5708e7b575b4b67;
      src125 <= 128'hc00276d8b6b3557b426d3948b4653341;
      src126 <= 128'h34f33a4ef835d15b4dbcf517e7c0dc23;
      src127 <= 128'h4f4aa95c35e98768a3a38fa5e8bf9cd8;
      #1
      src000 <= 128'h227b748ab4e2c460435b3a73d1cb8b27;
      src001 <= 128'h21a5123f38dd43bd3f97f4f8814c8efb;
      src002 <= 128'h5ccc0c1ddd5c4caf1a4e08cf7ee1f0e5;
      src003 <= 128'hb2564c0b219caedcb592fd3797a012e7;
      src004 <= 128'hebae29deb77920beddea624332d2f228;
      src005 <= 128'h9e34bd9b39f098da5bcdf979ed30655e;
      src006 <= 128'h523ac49a8a6a7ef20ac1f14676c8c182;
      src007 <= 128'h74af7dc29c4a8b3d71bd58f50b7865f;
      src008 <= 128'haa14625c39aa80fc2daa01238987a6fd;
      src009 <= 128'hb6608cf3b2e1d8481d87667a79b638c8;
      src010 <= 128'h9cec5333b416cbed01d580ec4a53ba16;
      src011 <= 128'h15f33777263c32210c099d16f195a9bb;
      src012 <= 128'hbacdd3134f9f9c7e41bc7237fff4f1fe;
      src013 <= 128'h9c16d57c968b1abdcef46fcc3954b25a;
      src014 <= 128'hf109bc67a0f80547d71388efc973c4e3;
      src015 <= 128'h30b3ede86b6d74ab2bb0e0065242b4a9;
      src016 <= 128'h8b3d5eb09aebda58c535693ef62bc9e4;
      src017 <= 128'hc5fd4007b2570a2e80746d98642d9ecc;
      src018 <= 128'h449c56ef3857ebe679ffa869834aac21;
      src019 <= 128'h9394eb115da6de86d849b508089711df;
      src020 <= 128'h90b89776cb77c423e5059533fa78c425;
      src021 <= 128'hb32c7f3c1cad91e87c36d70b60b9ad71;
      src022 <= 128'ha640d0f5f9eb611d327706c76ac04ece;
      src023 <= 128'h8abc0ff7c66e72f635dd3e7268fe2bdb;
      src024 <= 128'hbcab7a91183947ef579162f7d96be2f7;
      src025 <= 128'hea430e3ed5165c121af7f96ec0f9e07f;
      src026 <= 128'hf960229de1968f377781ea377ed8ce64;
      src027 <= 128'h9eef3cee5ef97498791d4347dd9fdc26;
      src028 <= 128'h910f8f667311274d0ca97ff3a2cfff86;
      src029 <= 128'h97bfe2e4f6df19473fff1ee0f5fddc69;
      src030 <= 128'h1c170895489594ed08dc3d4aad92540e;
      src031 <= 128'h5875de0f6a9000a8f74425c9563f4643;
      src032 <= 128'h20fc8e2974fb3857623fc5b9976d9953;
      src033 <= 128'h5fa8786e09bb66d83b2545c2287a302d;
      src034 <= 128'h4c2269c5b4d3669cbb65224f214140f5;
      src035 <= 128'h4ad99685861cd2f03206157cf5e32bfa;
      src036 <= 128'h1aa9210880d8241f4e4b41a12e21e8f7;
      src037 <= 128'hce0790d75f7e38982ddb2effdda72833;
      src038 <= 128'h632b16d24a14be4a41b1ea6a60e48300;
      src039 <= 128'hd252aac4f381331c95efbec5ef2d2a65;
      src040 <= 128'ha97e76efebefbae149c3a12df0bed3ed;
      src041 <= 128'hf0924ea87c837381958767902916bc05;
      src042 <= 128'he0dd1e208dfc0cb0dc97baec4fac816c;
      src043 <= 128'h4b86f79a7267eccc4e5a0edd7a1e3ce6;
      src044 <= 128'h763a98d72290b21334d2573b57db0c8b;
      src045 <= 128'h831520ca29d122e5e368fc63c94d1b10;
      src046 <= 128'h4e94228ca6107c6359245ab737c9f06d;
      src047 <= 128'h6eb7b98bb31190b621e4eb25adb2bb78;
      src048 <= 128'hf75f5cd55516c1a645d3fa2c08268550;
      src049 <= 128'h64426c12d8ea05db4c9ae79cb55dc17a;
      src050 <= 128'h9a4472e2de7ad23e2a0976e63faca756;
      src051 <= 128'hbca69710fcd3e74188ef1e2e73afe457;
      src052 <= 128'hd82c48259eb7e4e373df18f6484fca5f;
      src053 <= 128'h9295580eee6bf0de690aae3fade53235;
      src054 <= 128'h5cffd512e0309963114f17c1c4bd259f;
      src055 <= 128'h5962ceba2970243b3d47d3dfe97f9e57;
      src056 <= 128'h2c92f7725f779a39d619df9e7d1b254e;
      src057 <= 128'hd24a8ab9340794737edeb19d78020e02;
      src058 <= 128'hba4fa3cf84185d2d1ef4dec63a220bde;
      src059 <= 128'h39fd3acdd5b46772a4c7f528268ac0fc;
      src060 <= 128'h75af223a0f0ac1342e0d14ad8888d15e;
      src061 <= 128'h212589157b10077cbf32e5f786bbc79d;
      src062 <= 128'h99ac0892326e1c2f2fcfd8b73ceff664;
      src063 <= 128'h7b2846bac6c6e268597b322c572c55f1;
      src064 <= 128'h90a069ba5447353bc9dc6fb4f5677aaf;
      src065 <= 128'ha2af96924d735a4615dc9a2652b3fb34;
      src066 <= 128'hc7caa96bb098a39f12e903c1e33a8123;
      src067 <= 128'h412dfafafad63061ececa76bf30c85e;
      src068 <= 128'h8f484ea4144304640642485f3df629a3;
      src069 <= 128'h625237086d12f9cc4ea4f2ada8888536;
      src070 <= 128'hb9594d00f9cc2893b98857f8f098f6d8;
      src071 <= 128'h54496139add66d2053f3f048d814a978;
      src072 <= 128'hf654f453a5c23dc2cf8c01c4f23c7052;
      src073 <= 128'h6c7434eca59a476ccdcfefabe1f51fdc;
      src074 <= 128'h21c70fd7f4a9f3dc12cff12150909951;
      src075 <= 128'hb72cabfcf664107471f9d5190bd89c73;
      src076 <= 128'he675e7e7f848f19ad1fa1e143cde8704;
      src077 <= 128'hf9405ecf8c0f1c3e6aab5919a2cd8317;
      src078 <= 128'h9eabc602d98dee37e78297aacfd9a1d0;
      src079 <= 128'hf3e77c602cd395ebc2907413dcb2c15c;
      src080 <= 128'h3127f05b0a964cb9a62a24d01047111a;
      src081 <= 128'hcb562026a4d69d945097be87168d8bf9;
      src082 <= 128'hd54f5bd536ff84c82c7ce621f617ff9;
      src083 <= 128'h2b754b26e244aca8cd4ca3a2093c656e;
      src084 <= 128'h48d798785a4a65b6f3f2bcac5f927b3b;
      src085 <= 128'hc11bd09f6d0e08d4a819b75174380926;
      src086 <= 128'h3e6e6845bc97d93afb5c8295a67db9d6;
      src087 <= 128'h275ab60d7b1eaff70476d9681803b6e7;
      src088 <= 128'hd0bd1c4921a3d1c5408ebd5e17425e7;
      src089 <= 128'hcdc16eaf416b3bd285bfb8e58119d8a5;
      src090 <= 128'h514ae2ef9ba8b8f16a6103634cb0ffb0;
      src091 <= 128'h20b293a9b83d667c7e57bf3c0461d287;
      src092 <= 128'h400a67fc35ca4006085698d7a91b2a6f;
      src093 <= 128'h4b98a7b58116466930ca8e21b6522437;
      src094 <= 128'h36b7e56b6b1c08c4e469f10892894e79;
      src095 <= 128'hb4a9ed2c0123ce86d598baa1ad8bfe6d;
      src096 <= 128'h368f215b56d8e9f38a73d02868a08ddb;
      src097 <= 128'hf23d695213122a21662cd634b10b8e0;
      src098 <= 128'ha76d4b32212178c70ce131dceecec051;
      src099 <= 128'hb92f22881c70a1b71c24bcf687e8b9a7;
      src100 <= 128'h7c8f8514e1939b89d39013af682e543;
      src101 <= 128'hce6fb966032778728ffe34c082597982;
      src102 <= 128'h70069215929b5ca4020e76f02a336ef6;
      src103 <= 128'he7326e1f64b21ca69938b9e782b22d43;
      src104 <= 128'h8cff3e991e8e2d522ab9c1851af0ed28;
      src105 <= 128'h9a240f2d0295156027e6311e794daba2;
      src106 <= 128'h42810d571e63e89a379e1ff84c07db5d;
      src107 <= 128'h74c6ff01e67383496fc7a8bd8e5c9abf;
      src108 <= 128'h645e83f96b0b97731b1abf6e6b6343c5;
      src109 <= 128'hb79cdee60547ae0311818f74addb5678;
      src110 <= 128'h347a5655b7f852c5336e33e25b608086;
      src111 <= 128'hdf6a19856ecb0b067dcc900ae689bad6;
      src112 <= 128'h2c464f3d119e1d1c04408df3200465b8;
      src113 <= 128'ha2d6d8c81c38b00d96b687fe99f3b2f0;
      src114 <= 128'h8a03a812bf505b6894d4d43ac2959368;
      src115 <= 128'h933cc2c7a78a25da23a4164941eae059;
      src116 <= 128'h7f6e05a600b35a929e0394e76f34ae62;
      src117 <= 128'hcabd877d48be9890da9f454686003bbc;
      src118 <= 128'hed5dc37361d8d152bb7144375cbb509a;
      src119 <= 128'hd56da186ba13ca529bba3d9bb939626a;
      src120 <= 128'ha64f5e71f4abf9d5a33f0524b3536dcb;
      src121 <= 128'ha0b0dea7560ba7be6a2496d81c3bc04f;
      src122 <= 128'hb56acae6f7fa36fc5587e3c5571532b3;
      src123 <= 128'h56e9ae4150011d9d259ac3245e94d303;
      src124 <= 128'h1ac45edb9be6a1c738820ff2656930b8;
      src125 <= 128'hc18f41d46ab92d9f2569b532370539b;
      src126 <= 128'hb1db0a78f2fd8e7a1ddf3199a03cf061;
      src127 <= 128'h555e45653a581614376305247cb9ca3e;
      #1
      src000 <= 128'h77dcf7b27d97613f433ca80a1b3c9c49;
      src001 <= 128'h45abd40367418726203da6391e0e2ffd;
      src002 <= 128'heded413bb43f355f2a9df500ff2abd86;
      src003 <= 128'h3ef1b23be15e787afb1ab1d26a2edd95;
      src004 <= 128'h2cbdb877544f06ddc0eea397d4a6e349;
      src005 <= 128'hc78ad66d4a9bfc00192edd37379c05da;
      src006 <= 128'hbb0250b377059fa856be7bee667c4de7;
      src007 <= 128'h7523fcc12a4e9db93e507e0f8f040c54;
      src008 <= 128'h440c4ed5c1a8ccc35c33da3094fc085b;
      src009 <= 128'h29db292a4bf637b49430715803cd6178;
      src010 <= 128'hdb627a3de37f656971899b9470b600c4;
      src011 <= 128'h1511a3f9c46e1738790b1990a428da2e;
      src012 <= 128'h6fd4d110b7dedde9ac26cf5b77082bdc;
      src013 <= 128'hfc14e5c1977d226020bdbe66468dc95e;
      src014 <= 128'h791dc0c47f1363754f4394338a4d266f;
      src015 <= 128'h4f22070ded39abe091539f8f503618d0;
      src016 <= 128'h70f498cd6cb008dcb00c15523f0bf534;
      src017 <= 128'h2da2bcd58a8ed273ece12e8b05cc70a1;
      src018 <= 128'ha82c84abef10e37fcba93005c4022537;
      src019 <= 128'h54b9fb20aedb5e9e8fa16d27d7fc0059;
      src020 <= 128'h284884a255e5c1d9b0364ad9ee5be9b9;
      src021 <= 128'h18ca01b52b5deb8a645d327b7b19062c;
      src022 <= 128'h35152cbaec4ff6abea07cfddee9cee1f;
      src023 <= 128'h517f6188e95ef6ab6757f6578e1c5e6;
      src024 <= 128'h146672ad4b9e091349e19b4d61c668ce;
      src025 <= 128'h795300f74a1393ab39b3c49db26c687c;
      src026 <= 128'h1c16dc39049e3af0ceb4d20e3d0d4b35;
      src027 <= 128'hcab4e61dd109e20a1a5bfffe0a09ac26;
      src028 <= 128'hd2865c0177f7ad194ee5ddf0d996f125;
      src029 <= 128'h496679f874655798aabc1f902de48434;
      src030 <= 128'h211312e12e99dffa903e36cf18f205bb;
      src031 <= 128'h480c762aec319b23c7ff1268f14bbea9;
      src032 <= 128'h118d4e31c8b92445119c1d81b2836ea;
      src033 <= 128'hb046463493a7468c10c15f57fed68dc1;
      src034 <= 128'he589d4bc6d6d14b17c771ff7a6d15070;
      src035 <= 128'hb4901da8af3e614041c9edfe2ba1c841;
      src036 <= 128'hf36ff7ce505749979916e08e3b51a890;
      src037 <= 128'hd6a3b56eaa784730992ced0d3db37b8;
      src038 <= 128'h7ec29b33ed5c684be273b6120cb6021e;
      src039 <= 128'hb66ec5b1919a8f4a6d6180619e63256a;
      src040 <= 128'h4a51de416ac85f42a9c0fdec6c25aad6;
      src041 <= 128'hb9527fba397ce787f01688e4b43bcab8;
      src042 <= 128'h531e9571092770d286c56c4579dd6e75;
      src043 <= 128'hffb2e1c5e8b463bfc7e02623c6fc2166;
      src044 <= 128'h1240c5fa87b8a1f9e00e7ef4de3b68b8;
      src045 <= 128'hbe72fa1e45ef60dbe37872462f3342b5;
      src046 <= 128'h6fcc8b274dadbfb008b4f16f30a407e9;
      src047 <= 128'hf19d09dd9bb6cafb82acaff5159ee507;
      src048 <= 128'haa9bb48d2134b4aabc8f167a04d6466e;
      src049 <= 128'h85cf70dfce7f88c7df171830174271de;
      src050 <= 128'h5fe5162e9a726e897531b0bf28714114;
      src051 <= 128'h21acdfefc6f2aace07ecafc15dab06c4;
      src052 <= 128'h2a236a88f66ae1d6e484a48ef8eaf989;
      src053 <= 128'h6919102b9d2b0c26787edf5e3b88f47d;
      src054 <= 128'he15100dfb36f6e304c05e70346a1faed;
      src055 <= 128'hdd618829ef78cdcd3d12928d5fceaae6;
      src056 <= 128'hf99d4c7767a84e192304deaeeaa42fb7;
      src057 <= 128'he60d2adad2c8ffade980e670c0773fe0;
      src058 <= 128'h4a4fa6a208e58a37aeb6eef8eef72f9e;
      src059 <= 128'heecb810375f31bf45e96c772358221cc;
      src060 <= 128'hc3e6e03c20c5716a876a516f3a5bdc38;
      src061 <= 128'hb6e1da1824d8b7fed00cf571ff3a4992;
      src062 <= 128'h21fb641b67018feb0a3db26e992ddd24;
      src063 <= 128'h7a3e128f36042f2c61e0967891bcb727;
      src064 <= 128'h8a6fe77386dd3b65673ba5c0c7405160;
      src065 <= 128'hde5a69cdab957917bd042c350962d28;
      src066 <= 128'hf62c38ed9d99eb49f01eb4dfb15fd5e8;
      src067 <= 128'hf867760a8b0cbeb53c1a1eb74d03697;
      src068 <= 128'hf170b8cc152705e5003d0a83e5ccaf94;
      src069 <= 128'h1d8a5b3a3512ccaf45856260c5dfdbb2;
      src070 <= 128'h3b10563a313890278c286cd46461d43b;
      src071 <= 128'h71ec94327bf1b37039d22d0466c0c7;
      src072 <= 128'h842645209be1b42f4f118ed83a08493c;
      src073 <= 128'h991cbb26c189fcb97c0910961770a506;
      src074 <= 128'hec31a254074fbe492c73746464022306;
      src075 <= 128'h647611e9347bdfff1276bb2e185f9658;
      src076 <= 128'hadc8b698c723092995c08df88032a324;
      src077 <= 128'ha523be6d538ceb94ad7b70fad3b9f176;
      src078 <= 128'hc55965e157326bfde5c5fb71a8c37f6a;
      src079 <= 128'h164e43959404fbf673d6192089ffc1b;
      src080 <= 128'haffb6b09467365a7d11b3ec42a3c0c48;
      src081 <= 128'h375c61ff2331b26275b19d44d4d28851;
      src082 <= 128'h450174c91558f8ff23bb5a0d38d7874f;
      src083 <= 128'h2456240a667e116585faeb3786c2462;
      src084 <= 128'h3f2630e3b3cb362259c21586320cd721;
      src085 <= 128'hdb47982941ee6cf104c2e32cea56fc9c;
      src086 <= 128'h703fe5910975308593019febea40451f;
      src087 <= 128'h94bad83ee3c6cbee5bc0c198fa39ff70;
      src088 <= 128'h6028562ff6e405cda753625ca092979e;
      src089 <= 128'h604e263e574b411a66cfd52f52b1791a;
      src090 <= 128'hc1b3c26325c1827df19f370b83271dd;
      src091 <= 128'h905d811c1beff1ff58ddd411f5d2148c;
      src092 <= 128'h8344866204a4211a40e1a7683cd17950;
      src093 <= 128'hbf3e777a85573355b5f22c1d509e7263;
      src094 <= 128'h5209308edf7a78a660f65ad08a8f4951;
      src095 <= 128'hb326ca45892af03ba5adf53b3bc3373b;
      src096 <= 128'h15e00003d84d858b475b4c14f8462054;
      src097 <= 128'hddb2f3dae95528be759bf9c4d625e7c4;
      src098 <= 128'h36771ea6418b6d331551de12d856bbb0;
      src099 <= 128'h8ca9db0b53475d8a44baf4271e49dc9e;
      src100 <= 128'h271097f10f835c81fa55ad573f9cd6;
      src101 <= 128'h9907e4c01a254c4e7b21fb005c151b78;
      src102 <= 128'h43b545203b19e603aa0415586326ee35;
      src103 <= 128'h7bfed5c5d4c3aaaaeceb437aabbddadb;
      src104 <= 128'h6f7302d62bd99ae20726dd9e0738191;
      src105 <= 128'ha89a150dc26ff9f46c356df73a49cb04;
      src106 <= 128'h4f926225ad4f0f4917c1bb39cd66eb5d;
      src107 <= 128'h21ece55eb486af13cba51fd656793f06;
      src108 <= 128'h1a3afac9365c6e111cda0f4b1d749336;
      src109 <= 128'h315b14ae8017fb92320eed22b6e3e228;
      src110 <= 128'h3ce9f48b7ac4322ed8f8cb97b255814f;
      src111 <= 128'hc2bf07cbd2f4cf2e5887a3f19722dd1e;
      src112 <= 128'ha9f5e7b14e4bf176d87ae31a9673060a;
      src113 <= 128'h3541adbd131693967edd05ba2901cb3a;
      src114 <= 128'h9875f4f2bfd8130578cedc415cc93118;
      src115 <= 128'hf57458f9bd16b04f2cf6c298413b5c6d;
      src116 <= 128'ha637bc63dc4f6fb6dcd4ff33eede3c34;
      src117 <= 128'hcb4612010838d851ba231ecfa7a96066;
      src118 <= 128'hc7b2f3ea7c909c40e3ffb4bca2fa5a36;
      src119 <= 128'hca172bea9470a0ddd9990703398d034;
      src120 <= 128'h23e868bad3b2b82856d830a398c5c7d9;
      src121 <= 128'h5b5b1743ba9c3ff31f0d918f2662a1d2;
      src122 <= 128'h95a58f6f504e99a0dc07f7ba1aa1ad8f;
      src123 <= 128'he69fc01b5b8ea83740d4e357f3bbf976;
      src124 <= 128'h31a2baf81c660eb40e7cd3cf9067f465;
      src125 <= 128'h38af9fe5dd34d576507a69f617bab888;
      src126 <= 128'h8c47eae1859fe6378db5bc77341b6ada;
      src127 <= 128'h217546adb386ea067c1197462fe6c4ac;
   end
endmodule

