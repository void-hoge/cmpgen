module compressor(
      input wire [0:0] src000,
      input wire [1:0] src001,
      input wire [2:0] src002,
      input wire [3:0] src003,
      input wire [4:0] src004,
      input wire [5:0] src005,
      input wire [6:0] src006,
      input wire [7:0] src007,
      input wire [8:0] src008,
      input wire [9:0] src009,
      input wire [10:0] src010,
      input wire [11:0] src011,
      input wire [12:0] src012,
      input wire [13:0] src013,
      input wire [14:0] src014,
      input wire [15:0] src015,
      input wire [16:0] src016,
      input wire [17:0] src017,
      input wire [18:0] src018,
      input wire [19:0] src019,
      input wire [20:0] src020,
      input wire [21:0] src021,
      input wire [22:0] src022,
      input wire [23:0] src023,
      input wire [24:0] src024,
      input wire [25:0] src025,
      input wire [26:0] src026,
      input wire [27:0] src027,
      input wire [28:0] src028,
      input wire [29:0] src029,
      input wire [30:0] src030,
      input wire [31:0] src031,
      input wire [32:0] src032,
      input wire [33:0] src033,
      input wire [34:0] src034,
      input wire [35:0] src035,
      input wire [36:0] src036,
      input wire [37:0] src037,
      input wire [38:0] src038,
      input wire [39:0] src039,
      input wire [40:0] src040,
      input wire [41:0] src041,
      input wire [42:0] src042,
      input wire [43:0] src043,
      input wire [44:0] src044,
      input wire [45:0] src045,
      input wire [46:0] src046,
      input wire [47:0] src047,
      input wire [48:0] src048,
      input wire [49:0] src049,
      input wire [50:0] src050,
      input wire [51:0] src051,
      input wire [52:0] src052,
      input wire [53:0] src053,
      input wire [54:0] src054,
      input wire [55:0] src055,
      input wire [56:0] src056,
      input wire [57:0] src057,
      input wire [58:0] src058,
      input wire [59:0] src059,
      input wire [60:0] src060,
      input wire [61:0] src061,
      input wire [62:0] src062,
      input wire [63:0] src063,
      input wire [62:0] src064,
      input wire [61:0] src065,
      input wire [60:0] src066,
      input wire [59:0] src067,
      input wire [58:0] src068,
      input wire [57:0] src069,
      input wire [56:0] src070,
      input wire [55:0] src071,
      input wire [54:0] src072,
      input wire [53:0] src073,
      input wire [52:0] src074,
      input wire [51:0] src075,
      input wire [50:0] src076,
      input wire [49:0] src077,
      input wire [48:0] src078,
      input wire [47:0] src079,
      input wire [46:0] src080,
      input wire [45:0] src081,
      input wire [44:0] src082,
      input wire [43:0] src083,
      input wire [42:0] src084,
      input wire [41:0] src085,
      input wire [40:0] src086,
      input wire [39:0] src087,
      input wire [38:0] src088,
      input wire [37:0] src089,
      input wire [36:0] src090,
      input wire [35:0] src091,
      input wire [34:0] src092,
      input wire [33:0] src093,
      input wire [32:0] src094,
      input wire [31:0] src095,
      input wire [30:0] src096,
      input wire [29:0] src097,
      input wire [28:0] src098,
      input wire [27:0] src099,
      input wire [26:0] src100,
      input wire [25:0] src101,
      input wire [24:0] src102,
      input wire [23:0] src103,
      input wire [22:0] src104,
      input wire [21:0] src105,
      input wire [20:0] src106,
      input wire [19:0] src107,
      input wire [18:0] src108,
      input wire [17:0] src109,
      input wire [16:0] src110,
      input wire [15:0] src111,
      input wire [14:0] src112,
      input wire [13:0] src113,
      input wire [12:0] src114,
      input wire [11:0] src115,
      input wire [10:0] src116,
      input wire [9:0] src117,
      input wire [8:0] src118,
      input wire [7:0] src119,
      input wire [6:0] src120,
      input wire [5:0] src121,
      input wire [4:0] src122,
      input wire [3:0] src123,
      input wire [2:0] src124,
      input wire [1:0] src125,
      input wire [0:0] src126,
      output wire [0:0] dst000,
      output wire [0:0] dst001,
      output wire [0:0] dst002,
      output wire [0:0] dst003,
      output wire [0:0] dst004,
      output wire [1:0] dst005,
      output wire [1:0] dst006,
      output wire [0:0] dst007,
      output wire [0:0] dst008,
      output wire [1:0] dst009,
      output wire [1:0] dst010,
      output wire [1:0] dst011,
      output wire [0:0] dst012,
      output wire [1:0] dst013,
      output wire [1:0] dst014,
      output wire [1:0] dst015,
      output wire [1:0] dst016,
      output wire [1:0] dst017,
      output wire [1:0] dst018,
      output wire [1:0] dst019,
      output wire [1:0] dst020,
      output wire [0:0] dst021,
      output wire [1:0] dst022,
      output wire [1:0] dst023,
      output wire [0:0] dst024,
      output wire [1:0] dst025,
      output wire [1:0] dst026,
      output wire [1:0] dst027,
      output wire [1:0] dst028,
      output wire [1:0] dst029,
      output wire [1:0] dst030,
      output wire [1:0] dst031,
      output wire [1:0] dst032,
      output wire [1:0] dst033,
      output wire [1:0] dst034,
      output wire [1:0] dst035,
      output wire [0:0] dst036,
      output wire [1:0] dst037,
      output wire [1:0] dst038,
      output wire [1:0] dst039,
      output wire [1:0] dst040,
      output wire [1:0] dst041,
      output wire [1:0] dst042,
      output wire [1:0] dst043,
      output wire [1:0] dst044,
      output wire [1:0] dst045,
      output wire [1:0] dst046,
      output wire [1:0] dst047,
      output wire [1:0] dst048,
      output wire [1:0] dst049,
      output wire [1:0] dst050,
      output wire [1:0] dst051,
      output wire [1:0] dst052,
      output wire [1:0] dst053,
      output wire [1:0] dst054,
      output wire [1:0] dst055,
      output wire [1:0] dst056,
      output wire [1:0] dst057,
      output wire [1:0] dst058,
      output wire [1:0] dst059,
      output wire [1:0] dst060,
      output wire [1:0] dst061,
      output wire [1:0] dst062,
      output wire [1:0] dst063,
      output wire [1:0] dst064,
      output wire [1:0] dst065,
      output wire [1:0] dst066,
      output wire [1:0] dst067,
      output wire [1:0] dst068,
      output wire [1:0] dst069,
      output wire [1:0] dst070,
      output wire [1:0] dst071,
      output wire [1:0] dst072,
      output wire [1:0] dst073,
      output wire [1:0] dst074,
      output wire [1:0] dst075,
      output wire [1:0] dst076,
      output wire [1:0] dst077,
      output wire [1:0] dst078,
      output wire [1:0] dst079,
      output wire [1:0] dst080,
      output wire [1:0] dst081,
      output wire [1:0] dst082,
      output wire [1:0] dst083,
      output wire [1:0] dst084,
      output wire [1:0] dst085,
      output wire [1:0] dst086,
      output wire [1:0] dst087,
      output wire [1:0] dst088,
      output wire [1:0] dst089,
      output wire [1:0] dst090,
      output wire [1:0] dst091,
      output wire [1:0] dst092,
      output wire [1:0] dst093,
      output wire [1:0] dst094,
      output wire [1:0] dst095,
      output wire [1:0] dst096,
      output wire [1:0] dst097,
      output wire [1:0] dst098,
      output wire [1:0] dst099,
      output wire [1:0] dst100,
      output wire [1:0] dst101,
      output wire [1:0] dst102,
      output wire [1:0] dst103,
      output wire [1:0] dst104,
      output wire [1:0] dst105,
      output wire [1:0] dst106,
      output wire [1:0] dst107,
      output wire [1:0] dst108,
      output wire [1:0] dst109,
      output wire [1:0] dst110,
      output wire [1:0] dst111,
      output wire [1:0] dst112,
      output wire [1:0] dst113,
      output wire [1:0] dst114,
      output wire [0:0] dst115,
      output wire [1:0] dst116,
      output wire [1:0] dst117,
      output wire [1:0] dst118,
      output wire [1:0] dst119,
      output wire [1:0] dst120,
      output wire [1:0] dst121,
      output wire [0:0] dst122,
      output wire [0:0] dst123,
      output wire [1:0] dst124,
      output wire [1:0] dst125,
      output wire [0:0] dst126,
      output wire [1:0] dst127,
      output wire [0:0] dst128
   );
   wire [5:0] stage000;
   wire [6:0] stage001;
   wire [7:0] stage002;
   wire [11:0] stage003;
   wire [13:0] stage004;
   wire [30:0] stage005;
   wire [20:0] stage006;
   wire [34:0] stage007;
   wire [23:0] stage008;
   wire [44:0] stage009;
   wire [21:0] stage010;
   wire [38:0] stage011;
   wire [26:0] stage012;
   wire [38:0] stage013;
   wire [36:0] stage014;
   wire [41:0] stage015;
   wire [41:0] stage016;
   wire [64:0] stage017;
   wire [38:0] stage018;
   wire [55:0] stage019;
   wire [55:0] stage020;
   wire [49:0] stage021;
   wire [66:0] stage022;
   wire [64:0] stage023;
   wire [48:0] stage024;
   wire [69:0] stage025;
   wire [65:0] stage026;
   wire [97:0] stage027;
   wire [58:0] stage028;
   wire [69:0] stage029;
   wire [65:0] stage030;
   wire [73:0] stage031;
   wire [97:0] stage032;
   wire [58:0] stage033;
   wire [76:0] stage034;
   wire [72:0] stage035;
   wire [71:0] stage036;
   wire [78:0] stage037;
   wire [92:0] stage038;
   wire [73:0] stage039;
   wire [90:0] stage040;
   wire [87:0] stage041;
   wire [97:0] stage042;
   wire [92:0] stage043;
   wire [90:0] stage044;
   wire [90:0] stage045;
   wire [89:0] stage046;
   wire [113:0] stage047;
   wire [134:0] stage048;
   wire [101:0] stage049;
   wire [100:0] stage050;
   wire [87:0] stage051;
   wire [108:0] stage052;
   wire [139:0] stage053;
   wire [129:0] stage054;
   wire [123:0] stage055;
   wire [102:0] stage056;
   wire [99:0] stage057;
   wire [102:0] stage058;
   wire [117:0] stage059;
   wire [108:0] stage060;
   wire [136:0] stage061;
   wire [140:0] stage062;
   wire [145:0] stage063;
   wire [121:0] stage064;
   wire [129:0] stage065;
   wire [111:0] stage066;
   wire [124:0] stage067;
   wire [114:0] stage068;
   wire [123:0] stage069;
   wire [112:0] stage070;
   wire [119:0] stage071;
   wire [111:0] stage072;
   wire [102:0] stage073;
   wire [121:0] stage074;
   wire [100:0] stage075;
   wire [96:0] stage076;
   wire [103:0] stage077;
   wire [102:0] stage078;
   wire [120:0] stage079;
   wire [97:0] stage080;
   wire [102:0] stage081;
   wire [84:0] stage082;
   wire [89:0] stage083;
   wire [94:0] stage084;
   wire [89:0] stage085;
   wire [88:0] stage086;
   wire [76:0] stage087;
   wire [78:0] stage088;
   wire [83:0] stage089;
   wire [79:0] stage090;
   wire [88:0] stage091;
   wire [99:0] stage092;
   wire [93:0] stage093;
   wire [82:0] stage094;
   wire [88:0] stage095;
   wire [61:0] stage096;
   wire [69:0] stage097;
   wire [76:0] stage098;
   wire [55:0] stage099;
   wire [65:0] stage100;
   wire [51:0] stage101;
   wire [73:0] stage102;
   wire [59:0] stage103;
   wire [40:0] stage104;
   wire [81:0] stage105;
   wire [60:0] stage106;
   wire [37:0] stage107;
   wire [54:0] stage108;
   wire [38:0] stage109;
   wire [36:0] stage110;
   wire [48:0] stage111;
   wire [34:0] stage112;
   wire [45:0] stage113;
   wire [32:0] stage114;
   wire [48:0] stage115;
   wire [42:0] stage116;
   wire [30:0] stage117;
   wire [21:0] stage118;
   wire [29:0] stage119;
   wire [21:0] stage120;
   wire [21:0] stage121;
   wire [16:0] stage122;
   wire [15:0] stage123;
   wire [17:0] stage124;
   wire [11:0] stage125;
   wire [7:0] stage126;
   wire [3:0] stage127;
   wire [2:0] stage128;
   assign stage000[0:0] = src000;
   assign stage001[1:0] = src001;
   assign stage002[2:0] = src002;
   assign stage003[3:0] = src003;
   assign stage004[4:0] = src004;
   assign stage005[5:0] = src005;
   assign stage006[6:0] = src006;
   assign stage007[7:0] = src007;
   assign stage008[8:0] = src008;
   assign stage009[9:0] = src009;
   assign stage010[10:0] = src010;
   assign stage011[11:0] = src011;
   assign stage012[12:0] = src012;
   assign stage013[13:0] = src013;
   assign stage014[14:0] = src014;
   assign stage015[15:0] = src015;
   assign stage016[16:0] = src016;
   assign stage017[17:0] = src017;
   assign stage018[18:0] = src018;
   assign stage019[19:0] = src019;
   assign stage020[20:0] = src020;
   assign stage021[21:0] = src021;
   assign stage022[22:0] = src022;
   assign stage023[23:0] = src023;
   assign stage024[24:0] = src024;
   assign stage025[25:0] = src025;
   assign stage026[26:0] = src026;
   assign stage027[27:0] = src027;
   assign stage028[28:0] = src028;
   assign stage029[29:0] = src029;
   assign stage030[30:0] = src030;
   assign stage031[31:0] = src031;
   assign stage032[32:0] = src032;
   assign stage033[33:0] = src033;
   assign stage034[34:0] = src034;
   assign stage035[35:0] = src035;
   assign stage036[36:0] = src036;
   assign stage037[37:0] = src037;
   assign stage038[38:0] = src038;
   assign stage039[39:0] = src039;
   assign stage040[40:0] = src040;
   assign stage041[41:0] = src041;
   assign stage042[42:0] = src042;
   assign stage043[43:0] = src043;
   assign stage044[44:0] = src044;
   assign stage045[45:0] = src045;
   assign stage046[46:0] = src046;
   assign stage047[47:0] = src047;
   assign stage048[48:0] = src048;
   assign stage049[49:0] = src049;
   assign stage050[50:0] = src050;
   assign stage051[51:0] = src051;
   assign stage052[52:0] = src052;
   assign stage053[53:0] = src053;
   assign stage054[54:0] = src054;
   assign stage055[55:0] = src055;
   assign stage056[56:0] = src056;
   assign stage057[57:0] = src057;
   assign stage058[58:0] = src058;
   assign stage059[59:0] = src059;
   assign stage060[60:0] = src060;
   assign stage061[61:0] = src061;
   assign stage062[62:0] = src062;
   assign stage063[63:0] = src063;
   assign stage064[62:0] = src064;
   assign stage065[61:0] = src065;
   assign stage066[60:0] = src066;
   assign stage067[59:0] = src067;
   assign stage068[58:0] = src068;
   assign stage069[57:0] = src069;
   assign stage070[56:0] = src070;
   assign stage071[55:0] = src071;
   assign stage072[54:0] = src072;
   assign stage073[53:0] = src073;
   assign stage074[52:0] = src074;
   assign stage075[51:0] = src075;
   assign stage076[50:0] = src076;
   assign stage077[49:0] = src077;
   assign stage078[48:0] = src078;
   assign stage079[47:0] = src079;
   assign stage080[46:0] = src080;
   assign stage081[45:0] = src081;
   assign stage082[44:0] = src082;
   assign stage083[43:0] = src083;
   assign stage084[42:0] = src084;
   assign stage085[41:0] = src085;
   assign stage086[40:0] = src086;
   assign stage087[39:0] = src087;
   assign stage088[38:0] = src088;
   assign stage089[37:0] = src089;
   assign stage090[36:0] = src090;
   assign stage091[35:0] = src091;
   assign stage092[34:0] = src092;
   assign stage093[33:0] = src093;
   assign stage094[32:0] = src094;
   assign stage095[31:0] = src095;
   assign stage096[30:0] = src096;
   assign stage097[29:0] = src097;
   assign stage098[28:0] = src098;
   assign stage099[27:0] = src099;
   assign stage100[26:0] = src100;
   assign stage101[25:0] = src101;
   assign stage102[24:0] = src102;
   assign stage103[23:0] = src103;
   assign stage104[22:0] = src104;
   assign stage105[21:0] = src105;
   assign stage106[20:0] = src106;
   assign stage107[19:0] = src107;
   assign stage108[18:0] = src108;
   assign stage109[17:0] = src109;
   assign stage110[16:0] = src110;
   assign stage111[15:0] = src111;
   assign stage112[14:0] = src112;
   assign stage113[13:0] = src113;
   assign stage114[12:0] = src114;
   assign stage115[11:0] = src115;
   assign stage116[10:0] = src116;
   assign stage117[9:0] = src117;
   assign stage118[8:0] = src118;
   assign stage119[7:0] = src119;
   assign stage120[6:0] = src120;
   assign stage121[5:0] = src121;
   assign stage122[4:0] = src122;
   assign stage123[3:0] = src123;
   assign stage124[2:0] = src124;
   assign stage125[1:0] = src125;
   assign stage126[0:0] = src126;
   assign dst000 = stage000[5:5];
   assign dst001 = stage001[6:6];
   assign dst002 = stage002[7:7];
   assign dst003 = stage003[11:11];
   assign dst004 = stage004[13:13];
   assign dst005 = stage005[30:29];
   assign dst006 = stage006[20:19];
   assign dst007 = stage007[34:34];
   assign dst008 = stage008[23:23];
   assign dst009 = stage009[44:43];
   assign dst010 = stage010[21:20];
   assign dst011 = stage011[38:37];
   assign dst012 = stage012[26:26];
   assign dst013 = stage013[38:37];
   assign dst014 = stage014[36:35];
   assign dst015 = stage015[41:40];
   assign dst016 = stage016[41:40];
   assign dst017 = stage017[64:63];
   assign dst018 = stage018[38:37];
   assign dst019 = stage019[55:54];
   assign dst020 = stage020[55:54];
   assign dst021 = stage021[49:49];
   assign dst022 = stage022[66:65];
   assign dst023 = stage023[64:63];
   assign dst024 = stage024[48:48];
   assign dst025 = stage025[69:68];
   assign dst026 = stage026[65:64];
   assign dst027 = stage027[97:96];
   assign dst028 = stage028[58:57];
   assign dst029 = stage029[69:68];
   assign dst030 = stage030[65:64];
   assign dst031 = stage031[73:72];
   assign dst032 = stage032[97:96];
   assign dst033 = stage033[58:57];
   assign dst034 = stage034[76:75];
   assign dst035 = stage035[72:71];
   assign dst036 = stage036[71:71];
   assign dst037 = stage037[78:77];
   assign dst038 = stage038[92:91];
   assign dst039 = stage039[73:72];
   assign dst040 = stage040[90:89];
   assign dst041 = stage041[87:86];
   assign dst042 = stage042[97:96];
   assign dst043 = stage043[92:91];
   assign dst044 = stage044[90:89];
   assign dst045 = stage045[90:89];
   assign dst046 = stage046[89:88];
   assign dst047 = stage047[113:112];
   assign dst048 = stage048[134:133];
   assign dst049 = stage049[101:100];
   assign dst050 = stage050[100:99];
   assign dst051 = stage051[87:86];
   assign dst052 = stage052[108:107];
   assign dst053 = stage053[139:138];
   assign dst054 = stage054[129:128];
   assign dst055 = stage055[123:122];
   assign dst056 = stage056[102:101];
   assign dst057 = stage057[99:98];
   assign dst058 = stage058[102:101];
   assign dst059 = stage059[117:116];
   assign dst060 = stage060[108:107];
   assign dst061 = stage061[136:135];
   assign dst062 = stage062[140:139];
   assign dst063 = stage063[145:144];
   assign dst064 = stage064[121:120];
   assign dst065 = stage065[129:128];
   assign dst066 = stage066[111:110];
   assign dst067 = stage067[124:123];
   assign dst068 = stage068[114:113];
   assign dst069 = stage069[123:122];
   assign dst070 = stage070[112:111];
   assign dst071 = stage071[119:118];
   assign dst072 = stage072[111:110];
   assign dst073 = stage073[102:101];
   assign dst074 = stage074[121:120];
   assign dst075 = stage075[100:99];
   assign dst076 = stage076[96:95];
   assign dst077 = stage077[103:102];
   assign dst078 = stage078[102:101];
   assign dst079 = stage079[120:119];
   assign dst080 = stage080[97:96];
   assign dst081 = stage081[102:101];
   assign dst082 = stage082[84:83];
   assign dst083 = stage083[89:88];
   assign dst084 = stage084[94:93];
   assign dst085 = stage085[89:88];
   assign dst086 = stage086[88:87];
   assign dst087 = stage087[76:75];
   assign dst088 = stage088[78:77];
   assign dst089 = stage089[83:82];
   assign dst090 = stage090[79:78];
   assign dst091 = stage091[88:87];
   assign dst092 = stage092[99:98];
   assign dst093 = stage093[93:92];
   assign dst094 = stage094[82:81];
   assign dst095 = stage095[88:87];
   assign dst096 = stage096[61:60];
   assign dst097 = stage097[69:68];
   assign dst098 = stage098[76:75];
   assign dst099 = stage099[55:54];
   assign dst100 = stage100[65:64];
   assign dst101 = stage101[51:50];
   assign dst102 = stage102[73:72];
   assign dst103 = stage103[59:58];
   assign dst104 = stage104[40:39];
   assign dst105 = stage105[81:80];
   assign dst106 = stage106[60:59];
   assign dst107 = stage107[37:36];
   assign dst108 = stage108[54:53];
   assign dst109 = stage109[38:37];
   assign dst110 = stage110[36:35];
   assign dst111 = stage111[48:47];
   assign dst112 = stage112[34:33];
   assign dst113 = stage113[45:44];
   assign dst114 = stage114[32:31];
   assign dst115 = stage115[48:48];
   assign dst116 = stage116[42:41];
   assign dst117 = stage117[30:29];
   assign dst118 = stage118[21:20];
   assign dst119 = stage119[29:28];
   assign dst120 = stage120[21:20];
   assign dst121 = stage121[21:20];
   assign dst122 = stage122[16:16];
   assign dst123 = stage123[15:15];
   assign dst124 = stage124[17:16];
   assign dst125 = stage125[11:10];
   assign dst126 = stage126[7:7];
   assign dst127 = stage127[3:2];
   assign dst128 = stage128[2:2];
   gpc1_1 gpc1_1_0(
      {stage000[0]},
      {stage000[1]}
   );
   gpc1343_5 gpc1343_5_1(
      {stage001[0], stage001[1], 1'h0},
      {stage002[0], stage002[1], stage002[2], 1'h0},
      {stage003[0], stage003[1], stage003[2]},
      {stage004[0]},
      {stage005[6], stage004[5], stage003[4], stage002[3], stage001[2]}
   );
   gpc1_1 gpc1_1_2(
      {stage003[3]},
      {stage003[5]}
   );
   gpc1_1 gpc1_1_3(
      {stage004[1]},
      {stage004[6]}
   );
   gpc1_1 gpc1_1_4(
      {stage004[2]},
      {stage004[7]}
   );
   gpc1_1 gpc1_1_5(
      {stage004[3]},
      {stage004[8]}
   );
   gpc1_1 gpc1_1_6(
      {stage004[4]},
      {stage004[9]}
   );
   gpc1_1 gpc1_1_7(
      {stage005[0]},
      {stage005[7]}
   );
   gpc1_1 gpc1_1_8(
      {stage005[1]},
      {stage005[8]}
   );
   gpc1_1 gpc1_1_9(
      {stage005[2]},
      {stage005[9]}
   );
   gpc1_1 gpc1_1_10(
      {stage005[3]},
      {stage005[10]}
   );
   gpc1_1 gpc1_1_11(
      {stage005[4]},
      {stage005[11]}
   );
   gpc1_1 gpc1_1_12(
      {stage005[5]},
      {stage005[12]}
   );
   gpc1_1 gpc1_1_13(
      {stage006[0]},
      {stage006[7]}
   );
   gpc1_1 gpc1_1_14(
      {stage006[1]},
      {stage006[8]}
   );
   gpc1_1 gpc1_1_15(
      {stage006[2]},
      {stage006[9]}
   );
   gpc1_1 gpc1_1_16(
      {stage006[3]},
      {stage006[10]}
   );
   gpc1_1 gpc1_1_17(
      {stage006[4]},
      {stage006[11]}
   );
   gpc1_1 gpc1_1_18(
      {stage006[5]},
      {stage006[12]}
   );
   gpc1_1 gpc1_1_19(
      {stage006[6]},
      {stage006[13]}
   );
   gpc1_1 gpc1_1_20(
      {stage007[0]},
      {stage007[8]}
   );
   gpc1_1 gpc1_1_21(
      {stage007[1]},
      {stage007[9]}
   );
   gpc1_1 gpc1_1_22(
      {stage007[2]},
      {stage007[10]}
   );
   gpc1_1 gpc1_1_23(
      {stage007[3]},
      {stage007[11]}
   );
   gpc1_1 gpc1_1_24(
      {stage007[4]},
      {stage007[12]}
   );
   gpc1_1 gpc1_1_25(
      {stage007[5]},
      {stage007[13]}
   );
   gpc1_1 gpc1_1_26(
      {stage007[6]},
      {stage007[14]}
   );
   gpc1_1 gpc1_1_27(
      {stage007[7]},
      {stage007[15]}
   );
   gpc1_1 gpc1_1_28(
      {stage008[0]},
      {stage008[9]}
   );
   gpc1_1 gpc1_1_29(
      {stage008[1]},
      {stage008[10]}
   );
   gpc1_1 gpc1_1_30(
      {stage008[2]},
      {stage008[11]}
   );
   gpc1_1 gpc1_1_31(
      {stage008[3]},
      {stage008[12]}
   );
   gpc615_5 gpc615_5_32(
      {stage008[4], stage008[5], stage008[6], stage008[7], stage008[8]},
      {stage009[0]},
      {stage010[0], stage010[1], stage010[2], stage010[3], stage010[4], stage010[5]},
      {stage012[13], stage011[12], stage010[11], stage009[10], stage008[13]}
   );
   gpc1_1 gpc1_1_33(
      {stage009[1]},
      {stage009[11]}
   );
   gpc1_1 gpc1_1_34(
      {stage009[2]},
      {stage009[12]}
   );
   gpc1_1 gpc1_1_35(
      {stage009[3]},
      {stage009[13]}
   );
   gpc1_1 gpc1_1_36(
      {stage009[4]},
      {stage009[14]}
   );
   gpc1_1 gpc1_1_37(
      {stage009[5]},
      {stage009[15]}
   );
   gpc1_1 gpc1_1_38(
      {stage009[6]},
      {stage009[16]}
   );
   gpc1_1 gpc1_1_39(
      {stage009[7]},
      {stage009[17]}
   );
   gpc1_1 gpc1_1_40(
      {stage009[8]},
      {stage009[18]}
   );
   gpc1_1 gpc1_1_41(
      {stage009[9]},
      {stage009[19]}
   );
   gpc615_5 gpc615_5_42(
      {stage010[6], stage010[7], stage010[8], stage010[9], stage010[10]},
      {stage011[0]},
      {stage012[0], stage012[1], stage012[2], stage012[3], stage012[4], stage012[5]},
      {stage014[15], stage013[14], stage012[14], stage011[13], stage010[12]}
   );
   gpc1_1 gpc1_1_43(
      {stage011[1]},
      {stage011[14]}
   );
   gpc1_1 gpc1_1_44(
      {stage011[2]},
      {stage011[15]}
   );
   gpc1_1 gpc1_1_45(
      {stage011[3]},
      {stage011[16]}
   );
   gpc1_1 gpc1_1_46(
      {stage011[4]},
      {stage011[17]}
   );
   gpc1_1 gpc1_1_47(
      {stage011[5]},
      {stage011[18]}
   );
   gpc1_1 gpc1_1_48(
      {stage011[6]},
      {stage011[19]}
   );
   gpc1_1 gpc1_1_49(
      {stage011[7]},
      {stage011[20]}
   );
   gpc1_1 gpc1_1_50(
      {stage011[8]},
      {stage011[21]}
   );
   gpc1_1 gpc1_1_51(
      {stage011[9]},
      {stage011[22]}
   );
   gpc1_1 gpc1_1_52(
      {stage011[10]},
      {stage011[23]}
   );
   gpc1_1 gpc1_1_53(
      {stage011[11]},
      {stage011[24]}
   );
   gpc1_1 gpc1_1_54(
      {stage012[6]},
      {stage012[15]}
   );
   gpc606_5 gpc606_5_55(
      {stage012[7], stage012[8], stage012[9], stage012[10], stage012[11], stage012[12]},
      {stage014[0], stage014[1], stage014[2], stage014[3], stage014[4], stage014[5]},
      {stage016[17], stage015[16], stage014[16], stage013[15], stage012[16]}
   );
   gpc1_1 gpc1_1_56(
      {stage013[0]},
      {stage013[16]}
   );
   gpc1_1 gpc1_1_57(
      {stage013[1]},
      {stage013[17]}
   );
   gpc1_1 gpc1_1_58(
      {stage013[2]},
      {stage013[18]}
   );
   gpc1_1 gpc1_1_59(
      {stage013[3]},
      {stage013[19]}
   );
   gpc1_1 gpc1_1_60(
      {stage013[4]},
      {stage013[20]}
   );
   gpc1_1 gpc1_1_61(
      {stage013[5]},
      {stage013[21]}
   );
   gpc1_1 gpc1_1_62(
      {stage013[6]},
      {stage013[22]}
   );
   gpc1_1 gpc1_1_63(
      {stage013[7]},
      {stage013[23]}
   );
   gpc1_1 gpc1_1_64(
      {stage013[8]},
      {stage013[24]}
   );
   gpc1325_5 gpc1325_5_65(
      {stage013[9], stage013[10], stage013[11], stage013[12], stage013[13]},
      {stage014[6], stage014[7]},
      {stage015[0], stage015[1], stage015[2]},
      {stage016[0]},
      {stage017[18], stage016[18], stage015[17], stage014[17], stage013[25]}
   );
   gpc1_1 gpc1_1_66(
      {stage014[8]},
      {stage014[18]}
   );
   gpc1_1 gpc1_1_67(
      {stage014[9]},
      {stage014[19]}
   );
   gpc615_5 gpc615_5_68(
      {stage014[10], stage014[11], stage014[12], stage014[13], stage014[14]},
      {stage015[3]},
      {stage016[1], stage016[2], stage016[3], stage016[4], stage016[5], stage016[6]},
      {stage018[19], stage017[19], stage016[19], stage015[18], stage014[20]}
   );
   gpc1_1 gpc1_1_69(
      {stage015[4]},
      {stage015[19]}
   );
   gpc1_1 gpc1_1_70(
      {stage015[5]},
      {stage015[20]}
   );
   gpc1_1 gpc1_1_71(
      {stage015[6]},
      {stage015[21]}
   );
   gpc1_1 gpc1_1_72(
      {stage015[7]},
      {stage015[22]}
   );
   gpc1_1 gpc1_1_73(
      {stage015[8]},
      {stage015[23]}
   );
   gpc1_1 gpc1_1_74(
      {stage015[9]},
      {stage015[24]}
   );
   gpc606_5 gpc606_5_75(
      {stage015[10], stage015[11], stage015[12], stage015[13], stage015[14], stage015[15]},
      {stage017[0], stage017[1], stage017[2], stage017[3], stage017[4], stage017[5]},
      {stage019[20], stage018[20], stage017[20], stage016[20], stage015[25]}
   );
   gpc1_1 gpc1_1_76(
      {stage016[7]},
      {stage016[21]}
   );
   gpc1_1 gpc1_1_77(
      {stage016[8]},
      {stage016[22]}
   );
   gpc1_1 gpc1_1_78(
      {stage016[9]},
      {stage016[23]}
   );
   gpc1_1 gpc1_1_79(
      {stage016[10]},
      {stage016[24]}
   );
   gpc606_5 gpc606_5_80(
      {stage016[11], stage016[12], stage016[13], stage016[14], stage016[15], stage016[16]},
      {stage018[0], stage018[1], stage018[2], stage018[3], stage018[4], stage018[5]},
      {stage020[21], stage019[21], stage018[21], stage017[21], stage016[25]}
   );
   gpc1_1 gpc1_1_81(
      {stage017[6]},
      {stage017[22]}
   );
   gpc1_1 gpc1_1_82(
      {stage017[7]},
      {stage017[23]}
   );
   gpc1_1 gpc1_1_83(
      {stage017[8]},
      {stage017[24]}
   );
   gpc1_1 gpc1_1_84(
      {stage017[9]},
      {stage017[25]}
   );
   gpc1_1 gpc1_1_85(
      {stage017[10]},
      {stage017[26]}
   );
   gpc1_1 gpc1_1_86(
      {stage017[11]},
      {stage017[27]}
   );
   gpc1_1 gpc1_1_87(
      {stage017[12]},
      {stage017[28]}
   );
   gpc1_1 gpc1_1_88(
      {stage017[13]},
      {stage017[29]}
   );
   gpc1_1 gpc1_1_89(
      {stage017[14]},
      {stage017[30]}
   );
   gpc1_1 gpc1_1_90(
      {stage017[15]},
      {stage017[31]}
   );
   gpc1_1 gpc1_1_91(
      {stage017[16]},
      {stage017[32]}
   );
   gpc1_1 gpc1_1_92(
      {stage017[17]},
      {stage017[33]}
   );
   gpc1_1 gpc1_1_93(
      {stage018[6]},
      {stage018[22]}
   );
   gpc606_5 gpc606_5_94(
      {stage018[7], stage018[8], stage018[9], stage018[10], stage018[11], stage018[12]},
      {stage020[0], stage020[1], stage020[2], stage020[3], stage020[4], stage020[5]},
      {stage022[23], stage021[22], stage020[22], stage019[22], stage018[23]}
   );
   gpc606_5 gpc606_5_95(
      {stage018[13], stage018[14], stage018[15], stage018[16], stage018[17], stage018[18]},
      {stage020[6], stage020[7], stage020[8], stage020[9], stage020[10], stage020[11]},
      {stage022[24], stage021[23], stage020[23], stage019[23], stage018[24]}
   );
   gpc1_1 gpc1_1_96(
      {stage019[0]},
      {stage019[24]}
   );
   gpc1_1 gpc1_1_97(
      {stage019[1]},
      {stage019[25]}
   );
   gpc1_1 gpc1_1_98(
      {stage019[2]},
      {stage019[26]}
   );
   gpc1_1 gpc1_1_99(
      {stage019[3]},
      {stage019[27]}
   );
   gpc1_1 gpc1_1_100(
      {stage019[4]},
      {stage019[28]}
   );
   gpc1_1 gpc1_1_101(
      {stage019[5]},
      {stage019[29]}
   );
   gpc1_1 gpc1_1_102(
      {stage019[6]},
      {stage019[30]}
   );
   gpc1_1 gpc1_1_103(
      {stage019[7]},
      {stage019[31]}
   );
   gpc606_5 gpc606_5_104(
      {stage019[8], stage019[9], stage019[10], stage019[11], stage019[12], stage019[13]},
      {stage021[0], stage021[1], stage021[2], stage021[3], stage021[4], stage021[5]},
      {stage023[24], stage022[25], stage021[24], stage020[24], stage019[32]}
   );
   gpc606_5 gpc606_5_105(
      {stage019[14], stage019[15], stage019[16], stage019[17], stage019[18], stage019[19]},
      {stage021[6], stage021[7], stage021[8], stage021[9], stage021[10], stage021[11]},
      {stage023[25], stage022[26], stage021[25], stage020[25], stage019[33]}
   );
   gpc1_1 gpc1_1_106(
      {stage020[12]},
      {stage020[26]}
   );
   gpc1_1 gpc1_1_107(
      {stage020[13]},
      {stage020[27]}
   );
   gpc1_1 gpc1_1_108(
      {stage020[14]},
      {stage020[28]}
   );
   gpc1_1 gpc1_1_109(
      {stage020[15]},
      {stage020[29]}
   );
   gpc1_1 gpc1_1_110(
      {stage020[16]},
      {stage020[30]}
   );
   gpc1_1 gpc1_1_111(
      {stage020[17]},
      {stage020[31]}
   );
   gpc1_1 gpc1_1_112(
      {stage020[18]},
      {stage020[32]}
   );
   gpc1_1 gpc1_1_113(
      {stage020[19]},
      {stage020[33]}
   );
   gpc1_1 gpc1_1_114(
      {stage020[20]},
      {stage020[34]}
   );
   gpc1_1 gpc1_1_115(
      {stage021[12]},
      {stage021[26]}
   );
   gpc1_1 gpc1_1_116(
      {stage021[13]},
      {stage021[27]}
   );
   gpc1_1 gpc1_1_117(
      {stage021[14]},
      {stage021[28]}
   );
   gpc1_1 gpc1_1_118(
      {stage021[15]},
      {stage021[29]}
   );
   gpc1_1 gpc1_1_119(
      {stage021[16]},
      {stage021[30]}
   );
   gpc615_5 gpc615_5_120(
      {stage021[17], stage021[18], stage021[19], stage021[20], stage021[21]},
      {stage022[0]},
      {stage023[0], stage023[1], stage023[2], stage023[3], stage023[4], stage023[5]},
      {stage025[26], stage024[25], stage023[26], stage022[27], stage021[31]}
   );
   gpc1_1 gpc1_1_121(
      {stage022[1]},
      {stage022[28]}
   );
   gpc1_1 gpc1_1_122(
      {stage022[2]},
      {stage022[29]}
   );
   gpc1_1 gpc1_1_123(
      {stage022[3]},
      {stage022[30]}
   );
   gpc1_1 gpc1_1_124(
      {stage022[4]},
      {stage022[31]}
   );
   gpc1_1 gpc1_1_125(
      {stage022[5]},
      {stage022[32]}
   );
   gpc1_1 gpc1_1_126(
      {stage022[6]},
      {stage022[33]}
   );
   gpc1_1 gpc1_1_127(
      {stage022[7]},
      {stage022[34]}
   );
   gpc1_1 gpc1_1_128(
      {stage022[8]},
      {stage022[35]}
   );
   gpc1_1 gpc1_1_129(
      {stage022[9]},
      {stage022[36]}
   );
   gpc1_1 gpc1_1_130(
      {stage022[10]},
      {stage022[37]}
   );
   gpc1_1 gpc1_1_131(
      {stage022[11]},
      {stage022[38]}
   );
   gpc1_1 gpc1_1_132(
      {stage022[12]},
      {stage022[39]}
   );
   gpc615_5 gpc615_5_133(
      {stage022[13], stage022[14], stage022[15], stage022[16], stage022[17]},
      {stage023[6]},
      {stage024[0], stage024[1], stage024[2], stage024[3], stage024[4], stage024[5]},
      {stage026[27], stage025[27], stage024[26], stage023[27], stage022[40]}
   );
   gpc215_4 gpc215_4_134(
      {stage022[18], stage022[19], stage022[20], stage022[21], stage022[22]},
      {stage023[7]},
      {stage024[6], stage024[7]},
      {stage025[28], stage024[27], stage023[28], stage022[41]}
   );
   gpc1_1 gpc1_1_135(
      {stage023[8]},
      {stage023[29]}
   );
   gpc1_1 gpc1_1_136(
      {stage023[9]},
      {stage023[30]}
   );
   gpc1_1 gpc1_1_137(
      {stage023[10]},
      {stage023[31]}
   );
   gpc1_1 gpc1_1_138(
      {stage023[11]},
      {stage023[32]}
   );
   gpc1_1 gpc1_1_139(
      {stage023[12]},
      {stage023[33]}
   );
   gpc1_1 gpc1_1_140(
      {stage023[13]},
      {stage023[34]}
   );
   gpc1_1 gpc1_1_141(
      {stage023[14]},
      {stage023[35]}
   );
   gpc1_1 gpc1_1_142(
      {stage023[15]},
      {stage023[36]}
   );
   gpc1_1 gpc1_1_143(
      {stage023[16]},
      {stage023[37]}
   );
   gpc1_1 gpc1_1_144(
      {stage023[17]},
      {stage023[38]}
   );
   gpc1_1 gpc1_1_145(
      {stage023[18]},
      {stage023[39]}
   );
   gpc1_1 gpc1_1_146(
      {stage023[19]},
      {stage023[40]}
   );
   gpc1_1 gpc1_1_147(
      {stage023[20]},
      {stage023[41]}
   );
   gpc1_1 gpc1_1_148(
      {stage023[21]},
      {stage023[42]}
   );
   gpc1_1 gpc1_1_149(
      {stage023[22]},
      {stage023[43]}
   );
   gpc1_1 gpc1_1_150(
      {stage023[23]},
      {stage023[44]}
   );
   gpc1_1 gpc1_1_151(
      {stage024[8]},
      {stage024[28]}
   );
   gpc606_5 gpc606_5_152(
      {stage024[9], stage024[10], stage024[11], stage024[12], stage024[13], stage024[14]},
      {stage026[0], stage026[1], stage026[2], stage026[3], stage026[4], stage026[5]},
      {stage028[29], stage027[28], stage026[28], stage025[29], stage024[29]}
   );
   gpc2135_5 gpc2135_5_153(
      {stage024[15], stage024[16], stage024[17], stage024[18], stage024[19]},
      {stage025[0], stage025[1], stage025[2]},
      {stage026[6]},
      {stage027[0], stage027[1]},
      {stage028[30], stage027[29], stage026[29], stage025[30], stage024[30]}
   );
   gpc2135_5 gpc2135_5_154(
      {stage024[20], stage024[21], stage024[22], stage024[23], stage024[24]},
      {stage025[3], stage025[4], stage025[5]},
      {stage026[7]},
      {stage027[2], stage027[3]},
      {stage028[31], stage027[30], stage026[30], stage025[31], stage024[31]}
   );
   gpc1_1 gpc1_1_155(
      {stage025[6]},
      {stage025[32]}
   );
   gpc1_1 gpc1_1_156(
      {stage025[7]},
      {stage025[33]}
   );
   gpc1_1 gpc1_1_157(
      {stage025[8]},
      {stage025[34]}
   );
   gpc1_1 gpc1_1_158(
      {stage025[9]},
      {stage025[35]}
   );
   gpc1_1 gpc1_1_159(
      {stage025[10]},
      {stage025[36]}
   );
   gpc1_1 gpc1_1_160(
      {stage025[11]},
      {stage025[37]}
   );
   gpc1_1 gpc1_1_161(
      {stage025[12]},
      {stage025[38]}
   );
   gpc1_1 gpc1_1_162(
      {stage025[13]},
      {stage025[39]}
   );
   gpc1_1 gpc1_1_163(
      {stage025[14]},
      {stage025[40]}
   );
   gpc1_1 gpc1_1_164(
      {stage025[15]},
      {stage025[41]}
   );
   gpc1_1 gpc1_1_165(
      {stage025[16]},
      {stage025[42]}
   );
   gpc1_1 gpc1_1_166(
      {stage025[17]},
      {stage025[43]}
   );
   gpc1_1 gpc1_1_167(
      {stage025[18]},
      {stage025[44]}
   );
   gpc1_1 gpc1_1_168(
      {stage025[19]},
      {stage025[45]}
   );
   gpc1_1 gpc1_1_169(
      {stage025[20]},
      {stage025[46]}
   );
   gpc135_4 gpc135_4_170(
      {stage025[21], stage025[22], stage025[23], stage025[24], stage025[25]},
      {stage026[8], stage026[9], stage026[10]},
      {stage027[4]},
      {stage028[32], stage027[31], stage026[31], stage025[47]}
   );
   gpc1_1 gpc1_1_171(
      {stage026[11]},
      {stage026[32]}
   );
   gpc1_1 gpc1_1_172(
      {stage026[12]},
      {stage026[33]}
   );
   gpc1_1 gpc1_1_173(
      {stage026[13]},
      {stage026[34]}
   );
   gpc1_1 gpc1_1_174(
      {stage026[14]},
      {stage026[35]}
   );
   gpc1_1 gpc1_1_175(
      {stage026[15]},
      {stage026[36]}
   );
   gpc1_1 gpc1_1_176(
      {stage026[16]},
      {stage026[37]}
   );
   gpc1_1 gpc1_1_177(
      {stage026[17]},
      {stage026[38]}
   );
   gpc1_1 gpc1_1_178(
      {stage026[18]},
      {stage026[39]}
   );
   gpc1_1 gpc1_1_179(
      {stage026[19]},
      {stage026[40]}
   );
   gpc1_1 gpc1_1_180(
      {stage026[20]},
      {stage026[41]}
   );
   gpc606_5 gpc606_5_181(
      {stage026[21], stage026[22], stage026[23], stage026[24], stage026[25], stage026[26]},
      {stage028[0], stage028[1], stage028[2], stage028[3], stage028[4], stage028[5]},
      {stage030[31], stage029[30], stage028[33], stage027[32], stage026[42]}
   );
   gpc1_1 gpc1_1_182(
      {stage027[5]},
      {stage027[33]}
   );
   gpc1_1 gpc1_1_183(
      {stage027[6]},
      {stage027[34]}
   );
   gpc1_1 gpc1_1_184(
      {stage027[7]},
      {stage027[35]}
   );
   gpc1_1 gpc1_1_185(
      {stage027[8]},
      {stage027[36]}
   );
   gpc1_1 gpc1_1_186(
      {stage027[9]},
      {stage027[37]}
   );
   gpc1_1 gpc1_1_187(
      {stage027[10]},
      {stage027[38]}
   );
   gpc1_1 gpc1_1_188(
      {stage027[11]},
      {stage027[39]}
   );
   gpc1_1 gpc1_1_189(
      {stage027[12]},
      {stage027[40]}
   );
   gpc1_1 gpc1_1_190(
      {stage027[13]},
      {stage027[41]}
   );
   gpc1_1 gpc1_1_191(
      {stage027[14]},
      {stage027[42]}
   );
   gpc1_1 gpc1_1_192(
      {stage027[15]},
      {stage027[43]}
   );
   gpc1_1 gpc1_1_193(
      {stage027[16]},
      {stage027[44]}
   );
   gpc1_1 gpc1_1_194(
      {stage027[17]},
      {stage027[45]}
   );
   gpc1_1 gpc1_1_195(
      {stage027[18]},
      {stage027[46]}
   );
   gpc1_1 gpc1_1_196(
      {stage027[19]},
      {stage027[47]}
   );
   gpc1_1 gpc1_1_197(
      {stage027[20]},
      {stage027[48]}
   );
   gpc1_1 gpc1_1_198(
      {stage027[21]},
      {stage027[49]}
   );
   gpc1_1 gpc1_1_199(
      {stage027[22]},
      {stage027[50]}
   );
   gpc615_5 gpc615_5_200(
      {stage027[23], stage027[24], stage027[25], stage027[26], stage027[27]},
      {stage028[6]},
      {stage029[0], stage029[1], stage029[2], stage029[3], stage029[4], stage029[5]},
      {stage031[32], stage030[32], stage029[31], stage028[34], stage027[51]}
   );
   gpc1_1 gpc1_1_201(
      {stage028[7]},
      {stage028[35]}
   );
   gpc1_1 gpc1_1_202(
      {stage028[8]},
      {stage028[36]}
   );
   gpc615_5 gpc615_5_203(
      {stage028[9], stage028[10], stage028[11], stage028[12], stage028[13]},
      {stage029[6]},
      {stage030[0], stage030[1], stage030[2], stage030[3], stage030[4], stage030[5]},
      {stage032[33], stage031[33], stage030[33], stage029[32], stage028[37]}
   );
   gpc615_5 gpc615_5_204(
      {stage028[14], stage028[15], stage028[16], stage028[17], stage028[18]},
      {stage029[7]},
      {stage030[6], stage030[7], stage030[8], stage030[9], stage030[10], stage030[11]},
      {stage032[34], stage031[34], stage030[34], stage029[33], stage028[38]}
   );
   gpc615_5 gpc615_5_205(
      {stage028[19], stage028[20], stage028[21], stage028[22], stage028[23]},
      {stage029[8]},
      {stage030[12], stage030[13], stage030[14], stage030[15], stage030[16], stage030[17]},
      {stage032[35], stage031[35], stage030[35], stage029[34], stage028[39]}
   );
   gpc2135_5 gpc2135_5_206(
      {stage028[24], stage028[25], stage028[26], stage028[27], stage028[28]},
      {stage029[9], stage029[10], stage029[11]},
      {stage030[18]},
      {stage031[0], stage031[1]},
      {stage032[36], stage031[36], stage030[36], stage029[35], stage028[40]}
   );
   gpc1_1 gpc1_1_207(
      {stage029[12]},
      {stage029[36]}
   );
   gpc1_1 gpc1_1_208(
      {stage029[13]},
      {stage029[37]}
   );
   gpc1_1 gpc1_1_209(
      {stage029[14]},
      {stage029[38]}
   );
   gpc1_1 gpc1_1_210(
      {stage029[15]},
      {stage029[39]}
   );
   gpc1_1 gpc1_1_211(
      {stage029[16]},
      {stage029[40]}
   );
   gpc1_1 gpc1_1_212(
      {stage029[17]},
      {stage029[41]}
   );
   gpc1_1 gpc1_1_213(
      {stage029[18]},
      {stage029[42]}
   );
   gpc1_1 gpc1_1_214(
      {stage029[19]},
      {stage029[43]}
   );
   gpc1_1 gpc1_1_215(
      {stage029[20]},
      {stage029[44]}
   );
   gpc1_1 gpc1_1_216(
      {stage029[21]},
      {stage029[45]}
   );
   gpc1_1 gpc1_1_217(
      {stage029[22]},
      {stage029[46]}
   );
   gpc1_1 gpc1_1_218(
      {stage029[23]},
      {stage029[47]}
   );
   gpc606_5 gpc606_5_219(
      {stage029[24], stage029[25], stage029[26], stage029[27], stage029[28], stage029[29]},
      {stage031[2], stage031[3], stage031[4], stage031[5], stage031[6], stage031[7]},
      {stage033[34], stage032[37], stage031[37], stage030[37], stage029[48]}
   );
   gpc1_1 gpc1_1_220(
      {stage030[19]},
      {stage030[38]}
   );
   gpc1_1 gpc1_1_221(
      {stage030[20]},
      {stage030[39]}
   );
   gpc1_1 gpc1_1_222(
      {stage030[21]},
      {stage030[40]}
   );
   gpc1_1 gpc1_1_223(
      {stage030[22]},
      {stage030[41]}
   );
   gpc1_1 gpc1_1_224(
      {stage030[23]},
      {stage030[42]}
   );
   gpc1_1 gpc1_1_225(
      {stage030[24]},
      {stage030[43]}
   );
   gpc1_1 gpc1_1_226(
      {stage030[25]},
      {stage030[44]}
   );
   gpc615_5 gpc615_5_227(
      {stage030[26], stage030[27], stage030[28], stage030[29], stage030[30]},
      {stage031[8]},
      {stage032[0], stage032[1], stage032[2], stage032[3], stage032[4], stage032[5]},
      {stage034[35], stage033[35], stage032[38], stage031[38], stage030[45]}
   );
   gpc1_1 gpc1_1_228(
      {stage031[9]},
      {stage031[39]}
   );
   gpc1_1 gpc1_1_229(
      {stage031[10]},
      {stage031[40]}
   );
   gpc1_1 gpc1_1_230(
      {stage031[11]},
      {stage031[41]}
   );
   gpc1_1 gpc1_1_231(
      {stage031[12]},
      {stage031[42]}
   );
   gpc1_1 gpc1_1_232(
      {stage031[13]},
      {stage031[43]}
   );
   gpc1_1 gpc1_1_233(
      {stage031[14]},
      {stage031[44]}
   );
   gpc1_1 gpc1_1_234(
      {stage031[15]},
      {stage031[45]}
   );
   gpc1_1 gpc1_1_235(
      {stage031[16]},
      {stage031[46]}
   );
   gpc615_5 gpc615_5_236(
      {stage031[17], stage031[18], stage031[19], stage031[20], stage031[21]},
      {stage032[6]},
      {stage033[0], stage033[1], stage033[2], stage033[3], stage033[4], stage033[5]},
      {stage035[36], stage034[36], stage033[36], stage032[39], stage031[47]}
   );
   gpc615_5 gpc615_5_237(
      {stage031[22], stage031[23], stage031[24], stage031[25], stage031[26]},
      {stage032[7]},
      {stage033[6], stage033[7], stage033[8], stage033[9], stage033[10], stage033[11]},
      {stage035[37], stage034[37], stage033[37], stage032[40], stage031[48]}
   );
   gpc615_5 gpc615_5_238(
      {stage031[27], stage031[28], stage031[29], stage031[30], stage031[31]},
      {stage032[8]},
      {stage033[12], stage033[13], stage033[14], stage033[15], stage033[16], stage033[17]},
      {stage035[38], stage034[38], stage033[38], stage032[41], stage031[49]}
   );
   gpc1_1 gpc1_1_239(
      {stage032[9]},
      {stage032[42]}
   );
   gpc1_1 gpc1_1_240(
      {stage032[10]},
      {stage032[43]}
   );
   gpc1_1 gpc1_1_241(
      {stage032[11]},
      {stage032[44]}
   );
   gpc1_1 gpc1_1_242(
      {stage032[12]},
      {stage032[45]}
   );
   gpc1_1 gpc1_1_243(
      {stage032[13]},
      {stage032[46]}
   );
   gpc1_1 gpc1_1_244(
      {stage032[14]},
      {stage032[47]}
   );
   gpc1_1 gpc1_1_245(
      {stage032[15]},
      {stage032[48]}
   );
   gpc1_1 gpc1_1_246(
      {stage032[16]},
      {stage032[49]}
   );
   gpc1_1 gpc1_1_247(
      {stage032[17]},
      {stage032[50]}
   );
   gpc1_1 gpc1_1_248(
      {stage032[18]},
      {stage032[51]}
   );
   gpc1_1 gpc1_1_249(
      {stage032[19]},
      {stage032[52]}
   );
   gpc1_1 gpc1_1_250(
      {stage032[20]},
      {stage032[53]}
   );
   gpc1_1 gpc1_1_251(
      {stage032[21]},
      {stage032[54]}
   );
   gpc1_1 gpc1_1_252(
      {stage032[22]},
      {stage032[55]}
   );
   gpc1_1 gpc1_1_253(
      {stage032[23]},
      {stage032[56]}
   );
   gpc1_1 gpc1_1_254(
      {stage032[24]},
      {stage032[57]}
   );
   gpc1_1 gpc1_1_255(
      {stage032[25]},
      {stage032[58]}
   );
   gpc1_1 gpc1_1_256(
      {stage032[26]},
      {stage032[59]}
   );
   gpc1_1 gpc1_1_257(
      {stage032[27]},
      {stage032[60]}
   );
   gpc1_1 gpc1_1_258(
      {stage032[28]},
      {stage032[61]}
   );
   gpc1_1 gpc1_1_259(
      {stage032[29]},
      {stage032[62]}
   );
   gpc1_1 gpc1_1_260(
      {stage032[30]},
      {stage032[63]}
   );
   gpc1_1 gpc1_1_261(
      {stage032[31]},
      {stage032[64]}
   );
   gpc1_1 gpc1_1_262(
      {stage032[32]},
      {stage032[65]}
   );
   gpc1_1 gpc1_1_263(
      {stage033[18]},
      {stage033[39]}
   );
   gpc615_5 gpc615_5_264(
      {stage033[19], stage033[20], stage033[21], stage033[22], stage033[23]},
      {stage034[0]},
      {stage035[0], stage035[1], stage035[2], stage035[3], stage035[4], stage035[5]},
      {stage037[38], stage036[37], stage035[39], stage034[39], stage033[40]}
   );
   gpc615_5 gpc615_5_265(
      {stage033[24], stage033[25], stage033[26], stage033[27], stage033[28]},
      {stage034[1]},
      {stage035[6], stage035[7], stage035[8], stage035[9], stage035[10], stage035[11]},
      {stage037[39], stage036[38], stage035[40], stage034[40], stage033[41]}
   );
   gpc615_5 gpc615_5_266(
      {stage033[29], stage033[30], stage033[31], stage033[32], stage033[33]},
      {stage034[2]},
      {stage035[12], stage035[13], stage035[14], stage035[15], stage035[16], stage035[17]},
      {stage037[40], stage036[39], stage035[41], stage034[41], stage033[42]}
   );
   gpc1_1 gpc1_1_267(
      {stage034[3]},
      {stage034[42]}
   );
   gpc1_1 gpc1_1_268(
      {stage034[4]},
      {stage034[43]}
   );
   gpc1_1 gpc1_1_269(
      {stage034[5]},
      {stage034[44]}
   );
   gpc1_1 gpc1_1_270(
      {stage034[6]},
      {stage034[45]}
   );
   gpc1_1 gpc1_1_271(
      {stage034[7]},
      {stage034[46]}
   );
   gpc1_1 gpc1_1_272(
      {stage034[8]},
      {stage034[47]}
   );
   gpc1_1 gpc1_1_273(
      {stage034[9]},
      {stage034[48]}
   );
   gpc1_1 gpc1_1_274(
      {stage034[10]},
      {stage034[49]}
   );
   gpc1_1 gpc1_1_275(
      {stage034[11]},
      {stage034[50]}
   );
   gpc1_1 gpc1_1_276(
      {stage034[12]},
      {stage034[51]}
   );
   gpc1_1 gpc1_1_277(
      {stage034[13]},
      {stage034[52]}
   );
   gpc1_1 gpc1_1_278(
      {stage034[14]},
      {stage034[53]}
   );
   gpc615_5 gpc615_5_279(
      {stage034[15], stage034[16], stage034[17], stage034[18], stage034[19]},
      {stage035[18]},
      {stage036[0], stage036[1], stage036[2], stage036[3], stage036[4], stage036[5]},
      {stage038[39], stage037[41], stage036[40], stage035[42], stage034[54]}
   );
   gpc615_5 gpc615_5_280(
      {stage034[20], stage034[21], stage034[22], stage034[23], stage034[24]},
      {stage035[19]},
      {stage036[6], stage036[7], stage036[8], stage036[9], stage036[10], stage036[11]},
      {stage038[40], stage037[42], stage036[41], stage035[43], stage034[55]}
   );
   gpc615_5 gpc615_5_281(
      {stage034[25], stage034[26], stage034[27], stage034[28], stage034[29]},
      {stage035[20]},
      {stage036[12], stage036[13], stage036[14], stage036[15], stage036[16], stage036[17]},
      {stage038[41], stage037[43], stage036[42], stage035[44], stage034[56]}
   );
   gpc615_5 gpc615_5_282(
      {stage034[30], stage034[31], stage034[32], stage034[33], stage034[34]},
      {stage035[21]},
      {stage036[18], stage036[19], stage036[20], stage036[21], stage036[22], stage036[23]},
      {stage038[42], stage037[44], stage036[43], stage035[45], stage034[57]}
   );
   gpc1_1 gpc1_1_283(
      {stage035[22]},
      {stage035[46]}
   );
   gpc1_1 gpc1_1_284(
      {stage035[23]},
      {stage035[47]}
   );
   gpc606_5 gpc606_5_285(
      {stage035[24], stage035[25], stage035[26], stage035[27], stage035[28], stage035[29]},
      {stage037[0], stage037[1], stage037[2], stage037[3], stage037[4], stage037[5]},
      {stage039[40], stage038[43], stage037[45], stage036[44], stage035[48]}
   );
   gpc606_5 gpc606_5_286(
      {stage035[30], stage035[31], stage035[32], stage035[33], stage035[34], stage035[35]},
      {stage037[6], stage037[7], stage037[8], stage037[9], stage037[10], stage037[11]},
      {stage039[41], stage038[44], stage037[46], stage036[45], stage035[49]}
   );
   gpc1_1 gpc1_1_287(
      {stage036[24]},
      {stage036[46]}
   );
   gpc606_5 gpc606_5_288(
      {stage036[25], stage036[26], stage036[27], stage036[28], stage036[29], stage036[30]},
      {stage038[0], stage038[1], stage038[2], stage038[3], stage038[4], stage038[5]},
      {stage040[41], stage039[42], stage038[45], stage037[47], stage036[47]}
   );
   gpc606_5 gpc606_5_289(
      {stage036[31], stage036[32], stage036[33], stage036[34], stage036[35], stage036[36]},
      {stage038[6], stage038[7], stage038[8], stage038[9], stage038[10], stage038[11]},
      {stage040[42], stage039[43], stage038[46], stage037[48], stage036[48]}
   );
   gpc1_1 gpc1_1_290(
      {stage037[12]},
      {stage037[49]}
   );
   gpc1_1 gpc1_1_291(
      {stage037[13]},
      {stage037[50]}
   );
   gpc606_5 gpc606_5_292(
      {stage037[14], stage037[15], stage037[16], stage037[17], stage037[18], stage037[19]},
      {stage039[0], stage039[1], stage039[2], stage039[3], stage039[4], stage039[5]},
      {stage041[42], stage040[43], stage039[44], stage038[47], stage037[51]}
   );
   gpc606_5 gpc606_5_293(
      {stage037[20], stage037[21], stage037[22], stage037[23], stage037[24], stage037[25]},
      {stage039[6], stage039[7], stage039[8], stage039[9], stage039[10], stage039[11]},
      {stage041[43], stage040[44], stage039[45], stage038[48], stage037[52]}
   );
   gpc606_5 gpc606_5_294(
      {stage037[26], stage037[27], stage037[28], stage037[29], stage037[30], stage037[31]},
      {stage039[12], stage039[13], stage039[14], stage039[15], stage039[16], stage039[17]},
      {stage041[44], stage040[45], stage039[46], stage038[49], stage037[53]}
   );
   gpc606_5 gpc606_5_295(
      {stage037[32], stage037[33], stage037[34], stage037[35], stage037[36], stage037[37]},
      {stage039[18], stage039[19], stage039[20], stage039[21], stage039[22], stage039[23]},
      {stage041[45], stage040[46], stage039[47], stage038[50], stage037[54]}
   );
   gpc1_1 gpc1_1_296(
      {stage038[12]},
      {stage038[51]}
   );
   gpc1_1 gpc1_1_297(
      {stage038[13]},
      {stage038[52]}
   );
   gpc1_1 gpc1_1_298(
      {stage038[14]},
      {stage038[53]}
   );
   gpc1_1 gpc1_1_299(
      {stage038[15]},
      {stage038[54]}
   );
   gpc1_1 gpc1_1_300(
      {stage038[16]},
      {stage038[55]}
   );
   gpc1_1 gpc1_1_301(
      {stage038[17]},
      {stage038[56]}
   );
   gpc1_1 gpc1_1_302(
      {stage038[18]},
      {stage038[57]}
   );
   gpc1_1 gpc1_1_303(
      {stage038[19]},
      {stage038[58]}
   );
   gpc1_1 gpc1_1_304(
      {stage038[20]},
      {stage038[59]}
   );
   gpc1_1 gpc1_1_305(
      {stage038[21]},
      {stage038[60]}
   );
   gpc606_5 gpc606_5_306(
      {stage038[22], stage038[23], stage038[24], stage038[25], stage038[26], stage038[27]},
      {stage040[0], stage040[1], stage040[2], stage040[3], stage040[4], stage040[5]},
      {stage042[43], stage041[46], stage040[47], stage039[48], stage038[61]}
   );
   gpc606_5 gpc606_5_307(
      {stage038[28], stage038[29], stage038[30], stage038[31], stage038[32], stage038[33]},
      {stage040[6], stage040[7], stage040[8], stage040[9], stage040[10], stage040[11]},
      {stage042[44], stage041[47], stage040[48], stage039[49], stage038[62]}
   );
   gpc615_5 gpc615_5_308(
      {stage038[34], stage038[35], stage038[36], stage038[37], stage038[38]},
      {stage039[24]},
      {stage040[12], stage040[13], stage040[14], stage040[15], stage040[16], stage040[17]},
      {stage042[45], stage041[48], stage040[49], stage039[50], stage038[63]}
   );
   gpc1_1 gpc1_1_309(
      {stage039[25]},
      {stage039[51]}
   );
   gpc1_1 gpc1_1_310(
      {stage039[26]},
      {stage039[52]}
   );
   gpc1_1 gpc1_1_311(
      {stage039[27]},
      {stage039[53]}
   );
   gpc606_5 gpc606_5_312(
      {stage039[28], stage039[29], stage039[30], stage039[31], stage039[32], stage039[33]},
      {stage041[0], stage041[1], stage041[2], stage041[3], stage041[4], stage041[5]},
      {stage043[44], stage042[46], stage041[49], stage040[50], stage039[54]}
   );
   gpc606_5 gpc606_5_313(
      {stage039[34], stage039[35], stage039[36], stage039[37], stage039[38], stage039[39]},
      {stage041[6], stage041[7], stage041[8], stage041[9], stage041[10], stage041[11]},
      {stage043[45], stage042[47], stage041[50], stage040[51], stage039[55]}
   );
   gpc606_5 gpc606_5_314(
      {stage040[18], stage040[19], stage040[20], stage040[21], stage040[22], stage040[23]},
      {stage042[0], stage042[1], stage042[2], stage042[3], stage042[4], stage042[5]},
      {stage044[45], stage043[46], stage042[48], stage041[51], stage040[52]}
   );
   gpc606_5 gpc606_5_315(
      {stage040[24], stage040[25], stage040[26], stage040[27], stage040[28], stage040[29]},
      {stage042[6], stage042[7], stage042[8], stage042[9], stage042[10], stage042[11]},
      {stage044[46], stage043[47], stage042[49], stage041[52], stage040[53]}
   );
   gpc606_5 gpc606_5_316(
      {stage040[30], stage040[31], stage040[32], stage040[33], stage040[34], stage040[35]},
      {stage042[12], stage042[13], stage042[14], stage042[15], stage042[16], stage042[17]},
      {stage044[47], stage043[48], stage042[50], stage041[53], stage040[54]}
   );
   gpc606_5 gpc606_5_317(
      {stage040[36], stage040[37], stage040[38], stage040[39], stage040[40], 1'h0},
      {stage042[18], stage042[19], stage042[20], stage042[21], stage042[22], stage042[23]},
      {stage044[48], stage043[49], stage042[51], stage041[54], stage040[55]}
   );
   gpc1_1 gpc1_1_318(
      {stage041[12]},
      {stage041[55]}
   );
   gpc1_1 gpc1_1_319(
      {stage041[13]},
      {stage041[56]}
   );
   gpc1_1 gpc1_1_320(
      {stage041[14]},
      {stage041[57]}
   );
   gpc606_5 gpc606_5_321(
      {stage041[15], stage041[16], stage041[17], stage041[18], stage041[19], stage041[20]},
      {stage043[0], stage043[1], stage043[2], stage043[3], stage043[4], stage043[5]},
      {stage045[46], stage044[49], stage043[50], stage042[52], stage041[58]}
   );
   gpc606_5 gpc606_5_322(
      {stage041[21], stage041[22], stage041[23], stage041[24], stage041[25], stage041[26]},
      {stage043[6], stage043[7], stage043[8], stage043[9], stage043[10], stage043[11]},
      {stage045[47], stage044[50], stage043[51], stage042[53], stage041[59]}
   );
   gpc2135_5 gpc2135_5_323(
      {stage041[27], stage041[28], stage041[29], stage041[30], stage041[31]},
      {stage042[24], stage042[25], stage042[26]},
      {stage043[12]},
      {stage044[0], stage044[1]},
      {stage045[48], stage044[51], stage043[52], stage042[54], stage041[60]}
   );
   gpc2135_5 gpc2135_5_324(
      {stage041[32], stage041[33], stage041[34], stage041[35], stage041[36]},
      {stage042[27], stage042[28], stage042[29]},
      {stage043[13]},
      {stage044[2], stage044[3]},
      {stage045[49], stage044[52], stage043[53], stage042[55], stage041[61]}
   );
   gpc2135_5 gpc2135_5_325(
      {stage041[37], stage041[38], stage041[39], stage041[40], stage041[41]},
      {stage042[30], stage042[31], stage042[32]},
      {stage043[14]},
      {stage044[4], stage044[5]},
      {stage045[50], stage044[53], stage043[54], stage042[56], stage041[62]}
   );
   gpc1_1 gpc1_1_326(
      {stage042[33]},
      {stage042[57]}
   );
   gpc1_1 gpc1_1_327(
      {stage042[34]},
      {stage042[58]}
   );
   gpc1_1 gpc1_1_328(
      {stage042[35]},
      {stage042[59]}
   );
   gpc1_1 gpc1_1_329(
      {stage042[36]},
      {stage042[60]}
   );
   gpc1_1 gpc1_1_330(
      {stage042[37]},
      {stage042[61]}
   );
   gpc1_1 gpc1_1_331(
      {stage042[38]},
      {stage042[62]}
   );
   gpc1_1 gpc1_1_332(
      {stage042[39]},
      {stage042[63]}
   );
   gpc1_1 gpc1_1_333(
      {stage042[40]},
      {stage042[64]}
   );
   gpc1_1 gpc1_1_334(
      {stage042[41]},
      {stage042[65]}
   );
   gpc1_1 gpc1_1_335(
      {stage042[42]},
      {stage042[66]}
   );
   gpc1_1 gpc1_1_336(
      {stage043[15]},
      {stage043[55]}
   );
   gpc1_1 gpc1_1_337(
      {stage043[16]},
      {stage043[56]}
   );
   gpc1_1 gpc1_1_338(
      {stage043[17]},
      {stage043[57]}
   );
   gpc1_1 gpc1_1_339(
      {stage043[18]},
      {stage043[58]}
   );
   gpc1_1 gpc1_1_340(
      {stage043[19]},
      {stage043[59]}
   );
   gpc606_5 gpc606_5_341(
      {stage043[20], stage043[21], stage043[22], stage043[23], stage043[24], stage043[25]},
      {stage045[0], stage045[1], stage045[2], stage045[3], stage045[4], stage045[5]},
      {stage047[48], stage046[47], stage045[51], stage044[54], stage043[60]}
   );
   gpc606_5 gpc606_5_342(
      {stage043[26], stage043[27], stage043[28], stage043[29], stage043[30], stage043[31]},
      {stage045[6], stage045[7], stage045[8], stage045[9], stage045[10], stage045[11]},
      {stage047[49], stage046[48], stage045[52], stage044[55], stage043[61]}
   );
   gpc606_5 gpc606_5_343(
      {stage043[32], stage043[33], stage043[34], stage043[35], stage043[36], stage043[37]},
      {stage045[12], stage045[13], stage045[14], stage045[15], stage045[16], stage045[17]},
      {stage047[50], stage046[49], stage045[53], stage044[56], stage043[62]}
   );
   gpc606_5 gpc606_5_344(
      {stage043[38], stage043[39], stage043[40], stage043[41], stage043[42], stage043[43]},
      {stage045[18], stage045[19], stage045[20], stage045[21], stage045[22], stage045[23]},
      {stage047[51], stage046[50], stage045[54], stage044[57], stage043[63]}
   );
   gpc1_1 gpc1_1_345(
      {stage044[6]},
      {stage044[58]}
   );
   gpc1_1 gpc1_1_346(
      {stage044[7]},
      {stage044[59]}
   );
   gpc1_1 gpc1_1_347(
      {stage044[8]},
      {stage044[60]}
   );
   gpc1_1 gpc1_1_348(
      {stage044[9]},
      {stage044[61]}
   );
   gpc1_1 gpc1_1_349(
      {stage044[10]},
      {stage044[62]}
   );
   gpc1_1 gpc1_1_350(
      {stage044[11]},
      {stage044[63]}
   );
   gpc1_1 gpc1_1_351(
      {stage044[12]},
      {stage044[64]}
   );
   gpc1_1 gpc1_1_352(
      {stage044[13]},
      {stage044[65]}
   );
   gpc1_1 gpc1_1_353(
      {stage044[14]},
      {stage044[66]}
   );
   gpc606_5 gpc606_5_354(
      {stage044[15], stage044[16], stage044[17], stage044[18], stage044[19], stage044[20]},
      {stage046[0], stage046[1], stage046[2], stage046[3], stage046[4], stage046[5]},
      {stage048[49], stage047[52], stage046[51], stage045[55], stage044[67]}
   );
   gpc606_5 gpc606_5_355(
      {stage044[21], stage044[22], stage044[23], stage044[24], stage044[25], stage044[26]},
      {stage046[6], stage046[7], stage046[8], stage046[9], stage046[10], stage046[11]},
      {stage048[50], stage047[53], stage046[52], stage045[56], stage044[68]}
   );
   gpc606_5 gpc606_5_356(
      {stage044[27], stage044[28], stage044[29], stage044[30], stage044[31], stage044[32]},
      {stage046[12], stage046[13], stage046[14], stage046[15], stage046[16], stage046[17]},
      {stage048[51], stage047[54], stage046[53], stage045[57], stage044[69]}
   );
   gpc606_5 gpc606_5_357(
      {stage044[33], stage044[34], stage044[35], stage044[36], stage044[37], stage044[38]},
      {stage046[18], stage046[19], stage046[20], stage046[21], stage046[22], stage046[23]},
      {stage048[52], stage047[55], stage046[54], stage045[58], stage044[70]}
   );
   gpc606_5 gpc606_5_358(
      {stage044[39], stage044[40], stage044[41], stage044[42], stage044[43], stage044[44]},
      {stage046[24], stage046[25], stage046[26], stage046[27], stage046[28], stage046[29]},
      {stage048[53], stage047[56], stage046[55], stage045[59], stage044[71]}
   );
   gpc1_1 gpc1_1_359(
      {stage045[24]},
      {stage045[60]}
   );
   gpc1_1 gpc1_1_360(
      {stage045[25]},
      {stage045[61]}
   );
   gpc1_1 gpc1_1_361(
      {stage045[26]},
      {stage045[62]}
   );
   gpc1_1 gpc1_1_362(
      {stage045[27]},
      {stage045[63]}
   );
   gpc1_1 gpc1_1_363(
      {stage045[28]},
      {stage045[64]}
   );
   gpc1_1 gpc1_1_364(
      {stage045[29]},
      {stage045[65]}
   );
   gpc606_5 gpc606_5_365(
      {stage045[30], stage045[31], stage045[32], stage045[33], stage045[34], stage045[35]},
      {stage047[0], stage047[1], stage047[2], stage047[3], stage047[4], stage047[5]},
      {stage049[50], stage048[54], stage047[57], stage046[56], stage045[66]}
   );
   gpc615_5 gpc615_5_366(
      {stage045[36], stage045[37], stage045[38], stage045[39], stage045[40]},
      {stage046[30]},
      {stage047[6], stage047[7], stage047[8], stage047[9], stage047[10], stage047[11]},
      {stage049[51], stage048[55], stage047[58], stage046[57], stage045[67]}
   );
   gpc2135_5 gpc2135_5_367(
      {stage045[41], stage045[42], stage045[43], stage045[44], stage045[45]},
      {stage046[31], stage046[32], stage046[33]},
      {stage047[12]},
      {stage048[0], stage048[1]},
      {stage049[52], stage048[56], stage047[59], stage046[58], stage045[68]}
   );
   gpc1_1 gpc1_1_368(
      {stage046[34]},
      {stage046[59]}
   );
   gpc1_1 gpc1_1_369(
      {stage046[35]},
      {stage046[60]}
   );
   gpc623_5 gpc623_5_370(
      {stage046[36], stage046[37], stage046[38]},
      {stage047[13], stage047[14]},
      {stage048[2], stage048[3], stage048[4], stage048[5], stage048[6], stage048[7]},
      {stage050[51], stage049[53], stage048[57], stage047[60], stage046[61]}
   );
   gpc623_5 gpc623_5_371(
      {stage046[39], stage046[40], stage046[41]},
      {stage047[15], stage047[16]},
      {stage048[8], stage048[9], stage048[10], stage048[11], stage048[12], stage048[13]},
      {stage050[52], stage049[54], stage048[58], stage047[61], stage046[62]}
   );
   gpc1325_5 gpc1325_5_372(
      {stage046[42], stage046[43], stage046[44], stage046[45], stage046[46]},
      {stage047[17], stage047[18]},
      {stage048[14], stage048[15], stage048[16]},
      {stage049[0]},
      {stage050[53], stage049[55], stage048[59], stage047[62], stage046[63]}
   );
   gpc1_1 gpc1_1_373(
      {stage047[19]},
      {stage047[63]}
   );
   gpc1_1 gpc1_1_374(
      {stage047[20]},
      {stage047[64]}
   );
   gpc1_1 gpc1_1_375(
      {stage047[21]},
      {stage047[65]}
   );
   gpc1_1 gpc1_1_376(
      {stage047[22]},
      {stage047[66]}
   );
   gpc1_1 gpc1_1_377(
      {stage047[23]},
      {stage047[67]}
   );
   gpc1_1 gpc1_1_378(
      {stage047[24]},
      {stage047[68]}
   );
   gpc1_1 gpc1_1_379(
      {stage047[25]},
      {stage047[69]}
   );
   gpc1_1 gpc1_1_380(
      {stage047[26]},
      {stage047[70]}
   );
   gpc1_1 gpc1_1_381(
      {stage047[27]},
      {stage047[71]}
   );
   gpc1_1 gpc1_1_382(
      {stage047[28]},
      {stage047[72]}
   );
   gpc1_1 gpc1_1_383(
      {stage047[29]},
      {stage047[73]}
   );
   gpc1_1 gpc1_1_384(
      {stage047[30]},
      {stage047[74]}
   );
   gpc1_1 gpc1_1_385(
      {stage047[31]},
      {stage047[75]}
   );
   gpc1_1 gpc1_1_386(
      {stage047[32]},
      {stage047[76]}
   );
   gpc1_1 gpc1_1_387(
      {stage047[33]},
      {stage047[77]}
   );
   gpc1_1 gpc1_1_388(
      {stage047[34]},
      {stage047[78]}
   );
   gpc1_1 gpc1_1_389(
      {stage047[35]},
      {stage047[79]}
   );
   gpc1_1 gpc1_1_390(
      {stage047[36]},
      {stage047[80]}
   );
   gpc1_1 gpc1_1_391(
      {stage047[37]},
      {stage047[81]}
   );
   gpc1_1 gpc1_1_392(
      {stage047[38]},
      {stage047[82]}
   );
   gpc1_1 gpc1_1_393(
      {stage047[39]},
      {stage047[83]}
   );
   gpc1_1 gpc1_1_394(
      {stage047[40]},
      {stage047[84]}
   );
   gpc1_1 gpc1_1_395(
      {stage047[41]},
      {stage047[85]}
   );
   gpc1_1 gpc1_1_396(
      {stage047[42]},
      {stage047[86]}
   );
   gpc1_1 gpc1_1_397(
      {stage047[43]},
      {stage047[87]}
   );
   gpc1_1 gpc1_1_398(
      {stage047[44]},
      {stage047[88]}
   );
   gpc1_1 gpc1_1_399(
      {stage047[45]},
      {stage047[89]}
   );
   gpc1_1 gpc1_1_400(
      {stage047[46]},
      {stage047[90]}
   );
   gpc1_1 gpc1_1_401(
      {stage047[47]},
      {stage047[91]}
   );
   gpc1_1 gpc1_1_402(
      {stage048[17]},
      {stage048[60]}
   );
   gpc1_1 gpc1_1_403(
      {stage048[18]},
      {stage048[61]}
   );
   gpc1_1 gpc1_1_404(
      {stage048[19]},
      {stage048[62]}
   );
   gpc1_1 gpc1_1_405(
      {stage048[20]},
      {stage048[63]}
   );
   gpc1_1 gpc1_1_406(
      {stage048[21]},
      {stage048[64]}
   );
   gpc1_1 gpc1_1_407(
      {stage048[22]},
      {stage048[65]}
   );
   gpc1_1 gpc1_1_408(
      {stage048[23]},
      {stage048[66]}
   );
   gpc1_1 gpc1_1_409(
      {stage048[24]},
      {stage048[67]}
   );
   gpc1_1 gpc1_1_410(
      {stage048[25]},
      {stage048[68]}
   );
   gpc1_1 gpc1_1_411(
      {stage048[26]},
      {stage048[69]}
   );
   gpc1_1 gpc1_1_412(
      {stage048[27]},
      {stage048[70]}
   );
   gpc1_1 gpc1_1_413(
      {stage048[28]},
      {stage048[71]}
   );
   gpc1_1 gpc1_1_414(
      {stage048[29]},
      {stage048[72]}
   );
   gpc1_1 gpc1_1_415(
      {stage048[30]},
      {stage048[73]}
   );
   gpc1_1 gpc1_1_416(
      {stage048[31]},
      {stage048[74]}
   );
   gpc1_1 gpc1_1_417(
      {stage048[32]},
      {stage048[75]}
   );
   gpc1_1 gpc1_1_418(
      {stage048[33]},
      {stage048[76]}
   );
   gpc1_1 gpc1_1_419(
      {stage048[34]},
      {stage048[77]}
   );
   gpc1_1 gpc1_1_420(
      {stage048[35]},
      {stage048[78]}
   );
   gpc1_1 gpc1_1_421(
      {stage048[36]},
      {stage048[79]}
   );
   gpc1_1 gpc1_1_422(
      {stage048[37]},
      {stage048[80]}
   );
   gpc1_1 gpc1_1_423(
      {stage048[38]},
      {stage048[81]}
   );
   gpc1_1 gpc1_1_424(
      {stage048[39]},
      {stage048[82]}
   );
   gpc1_1 gpc1_1_425(
      {stage048[40]},
      {stage048[83]}
   );
   gpc1_1 gpc1_1_426(
      {stage048[41]},
      {stage048[84]}
   );
   gpc1_1 gpc1_1_427(
      {stage048[42]},
      {stage048[85]}
   );
   gpc606_5 gpc606_5_428(
      {stage048[43], stage048[44], stage048[45], stage048[46], stage048[47], stage048[48]},
      {stage050[0], stage050[1], stage050[2], stage050[3], stage050[4], stage050[5]},
      {stage052[53], stage051[52], stage050[54], stage049[56], stage048[86]}
   );
   gpc1_1 gpc1_1_429(
      {stage049[1]},
      {stage049[57]}
   );
   gpc1_1 gpc1_1_430(
      {stage049[2]},
      {stage049[58]}
   );
   gpc1_1 gpc1_1_431(
      {stage049[3]},
      {stage049[59]}
   );
   gpc1_1 gpc1_1_432(
      {stage049[4]},
      {stage049[60]}
   );
   gpc1_1 gpc1_1_433(
      {stage049[5]},
      {stage049[61]}
   );
   gpc1_1 gpc1_1_434(
      {stage049[6]},
      {stage049[62]}
   );
   gpc1_1 gpc1_1_435(
      {stage049[7]},
      {stage049[63]}
   );
   gpc1_1 gpc1_1_436(
      {stage049[8]},
      {stage049[64]}
   );
   gpc606_5 gpc606_5_437(
      {stage049[9], stage049[10], stage049[11], stage049[12], stage049[13], stage049[14]},
      {stage051[0], stage051[1], stage051[2], stage051[3], stage051[4], stage051[5]},
      {stage053[54], stage052[54], stage051[53], stage050[55], stage049[65]}
   );
   gpc606_5 gpc606_5_438(
      {stage049[15], stage049[16], stage049[17], stage049[18], stage049[19], stage049[20]},
      {stage051[6], stage051[7], stage051[8], stage051[9], stage051[10], stage051[11]},
      {stage053[55], stage052[55], stage051[54], stage050[56], stage049[66]}
   );
   gpc606_5 gpc606_5_439(
      {stage049[21], stage049[22], stage049[23], stage049[24], stage049[25], stage049[26]},
      {stage051[12], stage051[13], stage051[14], stage051[15], stage051[16], stage051[17]},
      {stage053[56], stage052[56], stage051[55], stage050[57], stage049[67]}
   );
   gpc606_5 gpc606_5_440(
      {stage049[27], stage049[28], stage049[29], stage049[30], stage049[31], stage049[32]},
      {stage051[18], stage051[19], stage051[20], stage051[21], stage051[22], stage051[23]},
      {stage053[57], stage052[57], stage051[56], stage050[58], stage049[68]}
   );
   gpc606_5 gpc606_5_441(
      {stage049[33], stage049[34], stage049[35], stage049[36], stage049[37], stage049[38]},
      {stage051[24], stage051[25], stage051[26], stage051[27], stage051[28], stage051[29]},
      {stage053[58], stage052[58], stage051[57], stage050[59], stage049[69]}
   );
   gpc606_5 gpc606_5_442(
      {stage049[39], stage049[40], stage049[41], stage049[42], stage049[43], stage049[44]},
      {stage051[30], stage051[31], stage051[32], stage051[33], stage051[34], stage051[35]},
      {stage053[59], stage052[59], stage051[58], stage050[60], stage049[70]}
   );
   gpc615_5 gpc615_5_443(
      {stage049[45], stage049[46], stage049[47], stage049[48], stage049[49]},
      {stage050[6]},
      {stage051[36], stage051[37], stage051[38], stage051[39], stage051[40], stage051[41]},
      {stage053[60], stage052[60], stage051[59], stage050[61], stage049[71]}
   );
   gpc1_1 gpc1_1_444(
      {stage050[7]},
      {stage050[62]}
   );
   gpc1_1 gpc1_1_445(
      {stage050[8]},
      {stage050[63]}
   );
   gpc1_1 gpc1_1_446(
      {stage050[9]},
      {stage050[64]}
   );
   gpc1_1 gpc1_1_447(
      {stage050[10]},
      {stage050[65]}
   );
   gpc1_1 gpc1_1_448(
      {stage050[11]},
      {stage050[66]}
   );
   gpc1_1 gpc1_1_449(
      {stage050[12]},
      {stage050[67]}
   );
   gpc1_1 gpc1_1_450(
      {stage050[13]},
      {stage050[68]}
   );
   gpc1_1 gpc1_1_451(
      {stage050[14]},
      {stage050[69]}
   );
   gpc606_5 gpc606_5_452(
      {stage050[15], stage050[16], stage050[17], stage050[18], stage050[19], stage050[20]},
      {stage052[0], stage052[1], stage052[2], stage052[3], stage052[4], stage052[5]},
      {stage054[55], stage053[61], stage052[61], stage051[60], stage050[70]}
   );
   gpc606_5 gpc606_5_453(
      {stage050[21], stage050[22], stage050[23], stage050[24], stage050[25], stage050[26]},
      {stage052[6], stage052[7], stage052[8], stage052[9], stage052[10], stage052[11]},
      {stage054[56], stage053[62], stage052[62], stage051[61], stage050[71]}
   );
   gpc606_5 gpc606_5_454(
      {stage050[27], stage050[28], stage050[29], stage050[30], stage050[31], stage050[32]},
      {stage052[12], stage052[13], stage052[14], stage052[15], stage052[16], stage052[17]},
      {stage054[57], stage053[63], stage052[63], stage051[62], stage050[72]}
   );
   gpc606_5 gpc606_5_455(
      {stage050[33], stage050[34], stage050[35], stage050[36], stage050[37], stage050[38]},
      {stage052[18], stage052[19], stage052[20], stage052[21], stage052[22], stage052[23]},
      {stage054[58], stage053[64], stage052[64], stage051[63], stage050[73]}
   );
   gpc606_5 gpc606_5_456(
      {stage050[39], stage050[40], stage050[41], stage050[42], stage050[43], stage050[44]},
      {stage052[24], stage052[25], stage052[26], stage052[27], stage052[28], stage052[29]},
      {stage054[59], stage053[65], stage052[65], stage051[64], stage050[74]}
   );
   gpc606_5 gpc606_5_457(
      {stage050[45], stage050[46], stage050[47], stage050[48], stage050[49], stage050[50]},
      {stage052[30], stage052[31], stage052[32], stage052[33], stage052[34], stage052[35]},
      {stage054[60], stage053[66], stage052[66], stage051[65], stage050[75]}
   );
   gpc615_5 gpc615_5_458(
      {stage051[42], stage051[43], stage051[44], stage051[45], stage051[46]},
      {stage052[36]},
      {stage053[0], stage053[1], stage053[2], stage053[3], stage053[4], stage053[5]},
      {stage055[56], stage054[61], stage053[67], stage052[67], stage051[66]}
   );
   gpc615_5 gpc615_5_459(
      {stage051[47], stage051[48], stage051[49], stage051[50], stage051[51]},
      {stage052[37]},
      {stage053[6], stage053[7], stage053[8], stage053[9], stage053[10], stage053[11]},
      {stage055[57], stage054[62], stage053[68], stage052[68], stage051[67]}
   );
   gpc1_1 gpc1_1_460(
      {stage052[38]},
      {stage052[69]}
   );
   gpc1_1 gpc1_1_461(
      {stage052[39]},
      {stage052[70]}
   );
   gpc1_1 gpc1_1_462(
      {stage052[40]},
      {stage052[71]}
   );
   gpc1_1 gpc1_1_463(
      {stage052[41]},
      {stage052[72]}
   );
   gpc1_1 gpc1_1_464(
      {stage052[42]},
      {stage052[73]}
   );
   gpc1_1 gpc1_1_465(
      {stage052[43]},
      {stage052[74]}
   );
   gpc1_1 gpc1_1_466(
      {stage052[44]},
      {stage052[75]}
   );
   gpc1_1 gpc1_1_467(
      {stage052[45]},
      {stage052[76]}
   );
   gpc1_1 gpc1_1_468(
      {stage052[46]},
      {stage052[77]}
   );
   gpc1_1 gpc1_1_469(
      {stage052[47]},
      {stage052[78]}
   );
   gpc1_1 gpc1_1_470(
      {stage052[48]},
      {stage052[79]}
   );
   gpc1_1 gpc1_1_471(
      {stage052[49]},
      {stage052[80]}
   );
   gpc1_1 gpc1_1_472(
      {stage052[50]},
      {stage052[81]}
   );
   gpc1_1 gpc1_1_473(
      {stage052[51]},
      {stage052[82]}
   );
   gpc1_1 gpc1_1_474(
      {stage052[52]},
      {stage052[83]}
   );
   gpc1_1 gpc1_1_475(
      {stage053[12]},
      {stage053[69]}
   );
   gpc1_1 gpc1_1_476(
      {stage053[13]},
      {stage053[70]}
   );
   gpc1_1 gpc1_1_477(
      {stage053[14]},
      {stage053[71]}
   );
   gpc1_1 gpc1_1_478(
      {stage053[15]},
      {stage053[72]}
   );
   gpc1_1 gpc1_1_479(
      {stage053[16]},
      {stage053[73]}
   );
   gpc1_1 gpc1_1_480(
      {stage053[17]},
      {stage053[74]}
   );
   gpc1_1 gpc1_1_481(
      {stage053[18]},
      {stage053[75]}
   );
   gpc1_1 gpc1_1_482(
      {stage053[19]},
      {stage053[76]}
   );
   gpc1_1 gpc1_1_483(
      {stage053[20]},
      {stage053[77]}
   );
   gpc1_1 gpc1_1_484(
      {stage053[21]},
      {stage053[78]}
   );
   gpc1_1 gpc1_1_485(
      {stage053[22]},
      {stage053[79]}
   );
   gpc1_1 gpc1_1_486(
      {stage053[23]},
      {stage053[80]}
   );
   gpc1_1 gpc1_1_487(
      {stage053[24]},
      {stage053[81]}
   );
   gpc1_1 gpc1_1_488(
      {stage053[25]},
      {stage053[82]}
   );
   gpc1_1 gpc1_1_489(
      {stage053[26]},
      {stage053[83]}
   );
   gpc1_1 gpc1_1_490(
      {stage053[27]},
      {stage053[84]}
   );
   gpc1_1 gpc1_1_491(
      {stage053[28]},
      {stage053[85]}
   );
   gpc1_1 gpc1_1_492(
      {stage053[29]},
      {stage053[86]}
   );
   gpc1_1 gpc1_1_493(
      {stage053[30]},
      {stage053[87]}
   );
   gpc1_1 gpc1_1_494(
      {stage053[31]},
      {stage053[88]}
   );
   gpc1_1 gpc1_1_495(
      {stage053[32]},
      {stage053[89]}
   );
   gpc1_1 gpc1_1_496(
      {stage053[33]},
      {stage053[90]}
   );
   gpc1_1 gpc1_1_497(
      {stage053[34]},
      {stage053[91]}
   );
   gpc1_1 gpc1_1_498(
      {stage053[35]},
      {stage053[92]}
   );
   gpc1_1 gpc1_1_499(
      {stage053[36]},
      {stage053[93]}
   );
   gpc1_1 gpc1_1_500(
      {stage053[37]},
      {stage053[94]}
   );
   gpc1_1 gpc1_1_501(
      {stage053[38]},
      {stage053[95]}
   );
   gpc1_1 gpc1_1_502(
      {stage053[39]},
      {stage053[96]}
   );
   gpc1_1 gpc1_1_503(
      {stage053[40]},
      {stage053[97]}
   );
   gpc1_1 gpc1_1_504(
      {stage053[41]},
      {stage053[98]}
   );
   gpc606_5 gpc606_5_505(
      {stage053[42], stage053[43], stage053[44], stage053[45], stage053[46], stage053[47]},
      {stage055[0], stage055[1], stage055[2], stage055[3], stage055[4], stage055[5]},
      {stage057[58], stage056[57], stage055[58], stage054[63], stage053[99]}
   );
   gpc606_5 gpc606_5_506(
      {stage053[48], stage053[49], stage053[50], stage053[51], stage053[52], stage053[53]},
      {stage055[6], stage055[7], stage055[8], stage055[9], stage055[10], stage055[11]},
      {stage057[59], stage056[58], stage055[59], stage054[64], stage053[100]}
   );
   gpc1_1 gpc1_1_507(
      {stage054[0]},
      {stage054[65]}
   );
   gpc1_1 gpc1_1_508(
      {stage054[1]},
      {stage054[66]}
   );
   gpc1_1 gpc1_1_509(
      {stage054[2]},
      {stage054[67]}
   );
   gpc1_1 gpc1_1_510(
      {stage054[3]},
      {stage054[68]}
   );
   gpc1_1 gpc1_1_511(
      {stage054[4]},
      {stage054[69]}
   );
   gpc1_1 gpc1_1_512(
      {stage054[5]},
      {stage054[70]}
   );
   gpc1_1 gpc1_1_513(
      {stage054[6]},
      {stage054[71]}
   );
   gpc1_1 gpc1_1_514(
      {stage054[7]},
      {stage054[72]}
   );
   gpc1_1 gpc1_1_515(
      {stage054[8]},
      {stage054[73]}
   );
   gpc1_1 gpc1_1_516(
      {stage054[9]},
      {stage054[74]}
   );
   gpc1_1 gpc1_1_517(
      {stage054[10]},
      {stage054[75]}
   );
   gpc1_1 gpc1_1_518(
      {stage054[11]},
      {stage054[76]}
   );
   gpc1_1 gpc1_1_519(
      {stage054[12]},
      {stage054[77]}
   );
   gpc1_1 gpc1_1_520(
      {stage054[13]},
      {stage054[78]}
   );
   gpc1_1 gpc1_1_521(
      {stage054[14]},
      {stage054[79]}
   );
   gpc1_1 gpc1_1_522(
      {stage054[15]},
      {stage054[80]}
   );
   gpc1_1 gpc1_1_523(
      {stage054[16]},
      {stage054[81]}
   );
   gpc1_1 gpc1_1_524(
      {stage054[17]},
      {stage054[82]}
   );
   gpc1_1 gpc1_1_525(
      {stage054[18]},
      {stage054[83]}
   );
   gpc1_1 gpc1_1_526(
      {stage054[19]},
      {stage054[84]}
   );
   gpc1_1 gpc1_1_527(
      {stage054[20]},
      {stage054[85]}
   );
   gpc1_1 gpc1_1_528(
      {stage054[21]},
      {stage054[86]}
   );
   gpc1_1 gpc1_1_529(
      {stage054[22]},
      {stage054[87]}
   );
   gpc1_1 gpc1_1_530(
      {stage054[23]},
      {stage054[88]}
   );
   gpc1_1 gpc1_1_531(
      {stage054[24]},
      {stage054[89]}
   );
   gpc1_1 gpc1_1_532(
      {stage054[25]},
      {stage054[90]}
   );
   gpc1_1 gpc1_1_533(
      {stage054[26]},
      {stage054[91]}
   );
   gpc1_1 gpc1_1_534(
      {stage054[27]},
      {stage054[92]}
   );
   gpc1_1 gpc1_1_535(
      {stage054[28]},
      {stage054[93]}
   );
   gpc1_1 gpc1_1_536(
      {stage054[29]},
      {stage054[94]}
   );
   gpc1_1 gpc1_1_537(
      {stage054[30]},
      {stage054[95]}
   );
   gpc606_5 gpc606_5_538(
      {stage054[31], stage054[32], stage054[33], stage054[34], stage054[35], stage054[36]},
      {stage056[0], stage056[1], stage056[2], stage056[3], stage056[4], stage056[5]},
      {stage058[59], stage057[60], stage056[59], stage055[60], stage054[96]}
   );
   gpc606_5 gpc606_5_539(
      {stage054[37], stage054[38], stage054[39], stage054[40], stage054[41], stage054[42]},
      {stage056[6], stage056[7], stage056[8], stage056[9], stage056[10], stage056[11]},
      {stage058[60], stage057[61], stage056[60], stage055[61], stage054[97]}
   );
   gpc606_5 gpc606_5_540(
      {stage054[43], stage054[44], stage054[45], stage054[46], stage054[47], stage054[48]},
      {stage056[12], stage056[13], stage056[14], stage056[15], stage056[16], stage056[17]},
      {stage058[61], stage057[62], stage056[61], stage055[62], stage054[98]}
   );
   gpc606_5 gpc606_5_541(
      {stage054[49], stage054[50], stage054[51], stage054[52], stage054[53], stage054[54]},
      {stage056[18], stage056[19], stage056[20], stage056[21], stage056[22], stage056[23]},
      {stage058[62], stage057[63], stage056[62], stage055[63], stage054[99]}
   );
   gpc1_1 gpc1_1_542(
      {stage055[12]},
      {stage055[64]}
   );
   gpc1_1 gpc1_1_543(
      {stage055[13]},
      {stage055[65]}
   );
   gpc1_1 gpc1_1_544(
      {stage055[14]},
      {stage055[66]}
   );
   gpc1_1 gpc1_1_545(
      {stage055[15]},
      {stage055[67]}
   );
   gpc1_1 gpc1_1_546(
      {stage055[16]},
      {stage055[68]}
   );
   gpc1_1 gpc1_1_547(
      {stage055[17]},
      {stage055[69]}
   );
   gpc1_1 gpc1_1_548(
      {stage055[18]},
      {stage055[70]}
   );
   gpc1_1 gpc1_1_549(
      {stage055[19]},
      {stage055[71]}
   );
   gpc1_1 gpc1_1_550(
      {stage055[20]},
      {stage055[72]}
   );
   gpc1_1 gpc1_1_551(
      {stage055[21]},
      {stage055[73]}
   );
   gpc1_1 gpc1_1_552(
      {stage055[22]},
      {stage055[74]}
   );
   gpc1_1 gpc1_1_553(
      {stage055[23]},
      {stage055[75]}
   );
   gpc1_1 gpc1_1_554(
      {stage055[24]},
      {stage055[76]}
   );
   gpc1_1 gpc1_1_555(
      {stage055[25]},
      {stage055[77]}
   );
   gpc615_5 gpc615_5_556(
      {stage055[26], stage055[27], stage055[28], stage055[29], stage055[30]},
      {stage056[24]},
      {stage057[0], stage057[1], stage057[2], stage057[3], stage057[4], stage057[5]},
      {stage059[60], stage058[63], stage057[64], stage056[63], stage055[78]}
   );
   gpc615_5 gpc615_5_557(
      {stage055[31], stage055[32], stage055[33], stage055[34], stage055[35]},
      {stage056[25]},
      {stage057[6], stage057[7], stage057[8], stage057[9], stage057[10], stage057[11]},
      {stage059[61], stage058[64], stage057[65], stage056[64], stage055[79]}
   );
   gpc615_5 gpc615_5_558(
      {stage055[36], stage055[37], stage055[38], stage055[39], stage055[40]},
      {stage056[26]},
      {stage057[12], stage057[13], stage057[14], stage057[15], stage057[16], stage057[17]},
      {stage059[62], stage058[65], stage057[66], stage056[65], stage055[80]}
   );
   gpc615_5 gpc615_5_559(
      {stage055[41], stage055[42], stage055[43], stage055[44], stage055[45]},
      {stage056[27]},
      {stage057[18], stage057[19], stage057[20], stage057[21], stage057[22], stage057[23]},
      {stage059[63], stage058[66], stage057[67], stage056[66], stage055[81]}
   );
   gpc615_5 gpc615_5_560(
      {stage055[46], stage055[47], stage055[48], stage055[49], stage055[50]},
      {stage056[28]},
      {stage057[24], stage057[25], stage057[26], stage057[27], stage057[28], stage057[29]},
      {stage059[64], stage058[67], stage057[68], stage056[67], stage055[82]}
   );
   gpc615_5 gpc615_5_561(
      {stage055[51], stage055[52], stage055[53], stage055[54], stage055[55]},
      {stage056[29]},
      {stage057[30], stage057[31], stage057[32], stage057[33], stage057[34], stage057[35]},
      {stage059[65], stage058[68], stage057[69], stage056[68], stage055[83]}
   );
   gpc1_1 gpc1_1_562(
      {stage056[30]},
      {stage056[69]}
   );
   gpc606_5 gpc606_5_563(
      {stage056[31], stage056[32], stage056[33], stage056[34], stage056[35], stage056[36]},
      {stage058[0], stage058[1], stage058[2], stage058[3], stage058[4], stage058[5]},
      {stage060[61], stage059[66], stage058[69], stage057[70], stage056[70]}
   );
   gpc615_5 gpc615_5_564(
      {stage056[37], stage056[38], stage056[39], stage056[40], stage056[41]},
      {stage057[36]},
      {stage058[6], stage058[7], stage058[8], stage058[9], stage058[10], stage058[11]},
      {stage060[62], stage059[67], stage058[70], stage057[71], stage056[71]}
   );
   gpc615_5 gpc615_5_565(
      {stage056[42], stage056[43], stage056[44], stage056[45], stage056[46]},
      {stage057[37]},
      {stage058[12], stage058[13], stage058[14], stage058[15], stage058[16], stage058[17]},
      {stage060[63], stage059[68], stage058[71], stage057[72], stage056[72]}
   );
   gpc615_5 gpc615_5_566(
      {stage056[47], stage056[48], stage056[49], stage056[50], stage056[51]},
      {stage057[38]},
      {stage058[18], stage058[19], stage058[20], stage058[21], stage058[22], stage058[23]},
      {stage060[64], stage059[69], stage058[72], stage057[73], stage056[73]}
   );
   gpc615_5 gpc615_5_567(
      {stage056[52], stage056[53], stage056[54], stage056[55], stage056[56]},
      {stage057[39]},
      {stage058[24], stage058[25], stage058[26], stage058[27], stage058[28], stage058[29]},
      {stage060[65], stage059[70], stage058[73], stage057[74], stage056[74]}
   );
   gpc1_1 gpc1_1_568(
      {stage057[40]},
      {stage057[75]}
   );
   gpc606_5 gpc606_5_569(
      {stage057[41], stage057[42], stage057[43], stage057[44], stage057[45], stage057[46]},
      {stage059[0], stage059[1], stage059[2], stage059[3], stage059[4], stage059[5]},
      {stage061[62], stage060[66], stage059[71], stage058[74], stage057[76]}
   );
   gpc606_5 gpc606_5_570(
      {stage057[47], stage057[48], stage057[49], stage057[50], stage057[51], stage057[52]},
      {stage059[6], stage059[7], stage059[8], stage059[9], stage059[10], stage059[11]},
      {stage061[63], stage060[67], stage059[72], stage058[75], stage057[77]}
   );
   gpc615_5 gpc615_5_571(
      {stage057[53], stage057[54], stage057[55], stage057[56], stage057[57]},
      {stage058[30]},
      {stage059[12], stage059[13], stage059[14], stage059[15], stage059[16], stage059[17]},
      {stage061[64], stage060[68], stage059[73], stage058[76], stage057[78]}
   );
   gpc615_5 gpc615_5_572(
      {stage058[31], stage058[32], stage058[33], stage058[34], stage058[35]},
      {stage059[18]},
      {stage060[0], stage060[1], stage060[2], stage060[3], stage060[4], stage060[5]},
      {stage062[63], stage061[65], stage060[69], stage059[74], stage058[77]}
   );
   gpc615_5 gpc615_5_573(
      {stage058[36], stage058[37], stage058[38], stage058[39], stage058[40]},
      {stage059[19]},
      {stage060[6], stage060[7], stage060[8], stage060[9], stage060[10], stage060[11]},
      {stage062[64], stage061[66], stage060[70], stage059[75], stage058[78]}
   );
   gpc615_5 gpc615_5_574(
      {stage058[41], stage058[42], stage058[43], stage058[44], stage058[45]},
      {stage059[20]},
      {stage060[12], stage060[13], stage060[14], stage060[15], stage060[16], stage060[17]},
      {stage062[65], stage061[67], stage060[71], stage059[76], stage058[79]}
   );
   gpc615_5 gpc615_5_575(
      {stage058[46], stage058[47], stage058[48], stage058[49], stage058[50]},
      {stage059[21]},
      {stage060[18], stage060[19], stage060[20], stage060[21], stage060[22], stage060[23]},
      {stage062[66], stage061[68], stage060[72], stage059[77], stage058[80]}
   );
   gpc615_5 gpc615_5_576(
      {stage058[51], stage058[52], stage058[53], stage058[54], stage058[55]},
      {stage059[22]},
      {stage060[24], stage060[25], stage060[26], stage060[27], stage060[28], stage060[29]},
      {stage062[67], stage061[69], stage060[73], stage059[78], stage058[81]}
   );
   gpc615_5 gpc615_5_577(
      {stage058[56], stage058[57], stage058[58], 1'h0, 1'h0},
      {stage059[23]},
      {stage060[30], stage060[31], stage060[32], stage060[33], stage060[34], stage060[35]},
      {stage062[68], stage061[70], stage060[74], stage059[79], stage058[82]}
   );
   gpc1_1 gpc1_1_578(
      {stage059[24]},
      {stage059[80]}
   );
   gpc1_1 gpc1_1_579(
      {stage059[25]},
      {stage059[81]}
   );
   gpc1_1 gpc1_1_580(
      {stage059[26]},
      {stage059[82]}
   );
   gpc1_1 gpc1_1_581(
      {stage059[27]},
      {stage059[83]}
   );
   gpc1_1 gpc1_1_582(
      {stage059[28]},
      {stage059[84]}
   );
   gpc606_5 gpc606_5_583(
      {stage059[29], stage059[30], stage059[31], stage059[32], stage059[33], stage059[34]},
      {stage061[0], stage061[1], stage061[2], stage061[3], stage061[4], stage061[5]},
      {stage063[64], stage062[69], stage061[71], stage060[75], stage059[85]}
   );
   gpc615_5 gpc615_5_584(
      {stage059[35], stage059[36], stage059[37], stage059[38], stage059[39]},
      {stage060[36]},
      {stage061[6], stage061[7], stage061[8], stage061[9], stage061[10], stage061[11]},
      {stage063[65], stage062[70], stage061[72], stage060[76], stage059[86]}
   );
   gpc615_5 gpc615_5_585(
      {stage059[40], stage059[41], stage059[42], stage059[43], stage059[44]},
      {stage060[37]},
      {stage061[12], stage061[13], stage061[14], stage061[15], stage061[16], stage061[17]},
      {stage063[66], stage062[71], stage061[73], stage060[77], stage059[87]}
   );
   gpc615_5 gpc615_5_586(
      {stage059[45], stage059[46], stage059[47], stage059[48], stage059[49]},
      {stage060[38]},
      {stage061[18], stage061[19], stage061[20], stage061[21], stage061[22], stage061[23]},
      {stage063[67], stage062[72], stage061[74], stage060[78], stage059[88]}
   );
   gpc615_5 gpc615_5_587(
      {stage059[50], stage059[51], stage059[52], stage059[53], stage059[54]},
      {stage060[39]},
      {stage061[24], stage061[25], stage061[26], stage061[27], stage061[28], stage061[29]},
      {stage063[68], stage062[73], stage061[75], stage060[79], stage059[89]}
   );
   gpc615_5 gpc615_5_588(
      {stage059[55], stage059[56], stage059[57], stage059[58], stage059[59]},
      {stage060[40]},
      {stage061[30], stage061[31], stage061[32], stage061[33], stage061[34], stage061[35]},
      {stage063[69], stage062[74], stage061[76], stage060[80], stage059[90]}
   );
   gpc615_5 gpc615_5_589(
      {stage060[41], stage060[42], stage060[43], stage060[44], stage060[45]},
      {stage061[36]},
      {stage062[0], stage062[1], stage062[2], stage062[3], stage062[4], stage062[5]},
      {stage064[63], stage063[70], stage062[75], stage061[77], stage060[81]}
   );
   gpc615_5 gpc615_5_590(
      {stage060[46], stage060[47], stage060[48], stage060[49], stage060[50]},
      {stage061[37]},
      {stage062[6], stage062[7], stage062[8], stage062[9], stage062[10], stage062[11]},
      {stage064[64], stage063[71], stage062[76], stage061[78], stage060[82]}
   );
   gpc615_5 gpc615_5_591(
      {stage060[51], stage060[52], stage060[53], stage060[54], stage060[55]},
      {stage061[38]},
      {stage062[12], stage062[13], stage062[14], stage062[15], stage062[16], stage062[17]},
      {stage064[65], stage063[72], stage062[77], stage061[79], stage060[83]}
   );
   gpc615_5 gpc615_5_592(
      {stage060[56], stage060[57], stage060[58], stage060[59], stage060[60]},
      {stage061[39]},
      {stage062[18], stage062[19], stage062[20], stage062[21], stage062[22], stage062[23]},
      {stage064[66], stage063[73], stage062[78], stage061[80], stage060[84]}
   );
   gpc1_1 gpc1_1_593(
      {stage061[40]},
      {stage061[81]}
   );
   gpc1_1 gpc1_1_594(
      {stage061[41]},
      {stage061[82]}
   );
   gpc1_1 gpc1_1_595(
      {stage061[42]},
      {stage061[83]}
   );
   gpc1_1 gpc1_1_596(
      {stage061[43]},
      {stage061[84]}
   );
   gpc1_1 gpc1_1_597(
      {stage061[44]},
      {stage061[85]}
   );
   gpc1_1 gpc1_1_598(
      {stage061[45]},
      {stage061[86]}
   );
   gpc1_1 gpc1_1_599(
      {stage061[46]},
      {stage061[87]}
   );
   gpc1_1 gpc1_1_600(
      {stage061[47]},
      {stage061[88]}
   );
   gpc1_1 gpc1_1_601(
      {stage061[48]},
      {stage061[89]}
   );
   gpc1_1 gpc1_1_602(
      {stage061[49]},
      {stage061[90]}
   );
   gpc1_1 gpc1_1_603(
      {stage061[50]},
      {stage061[91]}
   );
   gpc1_1 gpc1_1_604(
      {stage061[51]},
      {stage061[92]}
   );
   gpc1_1 gpc1_1_605(
      {stage061[52]},
      {stage061[93]}
   );
   gpc1_1 gpc1_1_606(
      {stage061[53]},
      {stage061[94]}
   );
   gpc1_1 gpc1_1_607(
      {stage061[54]},
      {stage061[95]}
   );
   gpc1_1 gpc1_1_608(
      {stage061[55]},
      {stage061[96]}
   );
   gpc1_1 gpc1_1_609(
      {stage061[56]},
      {stage061[97]}
   );
   gpc1_1 gpc1_1_610(
      {stage061[57]},
      {stage061[98]}
   );
   gpc1_1 gpc1_1_611(
      {stage061[58]},
      {stage061[99]}
   );
   gpc1_1 gpc1_1_612(
      {stage061[59]},
      {stage061[100]}
   );
   gpc1_1 gpc1_1_613(
      {stage061[60]},
      {stage061[101]}
   );
   gpc1_1 gpc1_1_614(
      {stage061[61]},
      {stage061[102]}
   );
   gpc1_1 gpc1_1_615(
      {stage062[24]},
      {stage062[79]}
   );
   gpc1_1 gpc1_1_616(
      {stage062[25]},
      {stage062[80]}
   );
   gpc1_1 gpc1_1_617(
      {stage062[26]},
      {stage062[81]}
   );
   gpc1_1 gpc1_1_618(
      {stage062[27]},
      {stage062[82]}
   );
   gpc1_1 gpc1_1_619(
      {stage062[28]},
      {stage062[83]}
   );
   gpc1_1 gpc1_1_620(
      {stage062[29]},
      {stage062[84]}
   );
   gpc1_1 gpc1_1_621(
      {stage062[30]},
      {stage062[85]}
   );
   gpc1_1 gpc1_1_622(
      {stage062[31]},
      {stage062[86]}
   );
   gpc1_1 gpc1_1_623(
      {stage062[32]},
      {stage062[87]}
   );
   gpc1_1 gpc1_1_624(
      {stage062[33]},
      {stage062[88]}
   );
   gpc1_1 gpc1_1_625(
      {stage062[34]},
      {stage062[89]}
   );
   gpc1_1 gpc1_1_626(
      {stage062[35]},
      {stage062[90]}
   );
   gpc1_1 gpc1_1_627(
      {stage062[36]},
      {stage062[91]}
   );
   gpc1_1 gpc1_1_628(
      {stage062[37]},
      {stage062[92]}
   );
   gpc1_1 gpc1_1_629(
      {stage062[38]},
      {stage062[93]}
   );
   gpc1_1 gpc1_1_630(
      {stage062[39]},
      {stage062[94]}
   );
   gpc1_1 gpc1_1_631(
      {stage062[40]},
      {stage062[95]}
   );
   gpc1_1 gpc1_1_632(
      {stage062[41]},
      {stage062[96]}
   );
   gpc1_1 gpc1_1_633(
      {stage062[42]},
      {stage062[97]}
   );
   gpc623_5 gpc623_5_634(
      {stage062[43], stage062[44], stage062[45]},
      {stage063[0], stage063[1]},
      {stage064[0], stage064[1], stage064[2], stage064[3], stage064[4], stage064[5]},
      {stage066[61], stage065[62], stage064[67], stage063[74], stage062[98]}
   );
   gpc606_5 gpc606_5_635(
      {stage062[46], stage062[47], stage062[48], stage062[49], stage062[50], stage062[51]},
      {stage064[6], stage064[7], stage064[8], stage064[9], stage064[10], stage064[11]},
      {stage066[62], stage065[63], stage064[68], stage063[75], stage062[99]}
   );
   gpc606_5 gpc606_5_636(
      {stage062[52], stage062[53], stage062[54], stage062[55], stage062[56], stage062[57]},
      {stage064[12], stage064[13], stage064[14], stage064[15], stage064[16], stage064[17]},
      {stage066[63], stage065[64], stage064[69], stage063[76], stage062[100]}
   );
   gpc615_5 gpc615_5_637(
      {stage062[58], stage062[59], stage062[60], stage062[61], stage062[62]},
      {stage063[2]},
      {stage064[18], stage064[19], stage064[20], stage064[21], stage064[22], stage064[23]},
      {stage066[64], stage065[65], stage064[70], stage063[77], stage062[101]}
   );
   gpc1_1 gpc1_1_638(
      {stage063[3]},
      {stage063[78]}
   );
   gpc1_1 gpc1_1_639(
      {stage063[4]},
      {stage063[79]}
   );
   gpc1_1 gpc1_1_640(
      {stage063[5]},
      {stage063[80]}
   );
   gpc1_1 gpc1_1_641(
      {stage063[6]},
      {stage063[81]}
   );
   gpc1_1 gpc1_1_642(
      {stage063[7]},
      {stage063[82]}
   );
   gpc1_1 gpc1_1_643(
      {stage063[8]},
      {stage063[83]}
   );
   gpc1_1 gpc1_1_644(
      {stage063[9]},
      {stage063[84]}
   );
   gpc1_1 gpc1_1_645(
      {stage063[10]},
      {stage063[85]}
   );
   gpc1_1 gpc1_1_646(
      {stage063[11]},
      {stage063[86]}
   );
   gpc1_1 gpc1_1_647(
      {stage063[12]},
      {stage063[87]}
   );
   gpc1_1 gpc1_1_648(
      {stage063[13]},
      {stage063[88]}
   );
   gpc1_1 gpc1_1_649(
      {stage063[14]},
      {stage063[89]}
   );
   gpc1_1 gpc1_1_650(
      {stage063[15]},
      {stage063[90]}
   );
   gpc1_1 gpc1_1_651(
      {stage063[16]},
      {stage063[91]}
   );
   gpc1_1 gpc1_1_652(
      {stage063[17]},
      {stage063[92]}
   );
   gpc1_1 gpc1_1_653(
      {stage063[18]},
      {stage063[93]}
   );
   gpc1_1 gpc1_1_654(
      {stage063[19]},
      {stage063[94]}
   );
   gpc1_1 gpc1_1_655(
      {stage063[20]},
      {stage063[95]}
   );
   gpc1_1 gpc1_1_656(
      {stage063[21]},
      {stage063[96]}
   );
   gpc606_5 gpc606_5_657(
      {stage063[22], stage063[23], stage063[24], stage063[25], stage063[26], stage063[27]},
      {stage065[0], stage065[1], stage065[2], stage065[3], stage065[4], stage065[5]},
      {stage067[60], stage066[65], stage065[66], stage064[71], stage063[97]}
   );
   gpc606_5 gpc606_5_658(
      {stage063[28], stage063[29], stage063[30], stage063[31], stage063[32], stage063[33]},
      {stage065[6], stage065[7], stage065[8], stage065[9], stage065[10], stage065[11]},
      {stage067[61], stage066[66], stage065[67], stage064[72], stage063[98]}
   );
   gpc606_5 gpc606_5_659(
      {stage063[34], stage063[35], stage063[36], stage063[37], stage063[38], stage063[39]},
      {stage065[12], stage065[13], stage065[14], stage065[15], stage065[16], stage065[17]},
      {stage067[62], stage066[67], stage065[68], stage064[73], stage063[99]}
   );
   gpc606_5 gpc606_5_660(
      {stage063[40], stage063[41], stage063[42], stage063[43], stage063[44], stage063[45]},
      {stage065[18], stage065[19], stage065[20], stage065[21], stage065[22], stage065[23]},
      {stage067[63], stage066[68], stage065[69], stage064[74], stage063[100]}
   );
   gpc606_5 gpc606_5_661(
      {stage063[46], stage063[47], stage063[48], stage063[49], stage063[50], stage063[51]},
      {stage065[24], stage065[25], stage065[26], stage065[27], stage065[28], stage065[29]},
      {stage067[64], stage066[69], stage065[70], stage064[75], stage063[101]}
   );
   gpc606_5 gpc606_5_662(
      {stage063[52], stage063[53], stage063[54], stage063[55], stage063[56], stage063[57]},
      {stage065[30], stage065[31], stage065[32], stage065[33], stage065[34], stage065[35]},
      {stage067[65], stage066[70], stage065[71], stage064[76], stage063[102]}
   );
   gpc606_5 gpc606_5_663(
      {stage063[58], stage063[59], stage063[60], stage063[61], stage063[62], stage063[63]},
      {stage065[36], stage065[37], stage065[38], stage065[39], stage065[40], stage065[41]},
      {stage067[66], stage066[71], stage065[72], stage064[77], stage063[103]}
   );
   gpc1_1 gpc1_1_664(
      {stage064[24]},
      {stage064[78]}
   );
   gpc1_1 gpc1_1_665(
      {stage064[25]},
      {stage064[79]}
   );
   gpc1_1 gpc1_1_666(
      {stage064[26]},
      {stage064[80]}
   );
   gpc1_1 gpc1_1_667(
      {stage064[27]},
      {stage064[81]}
   );
   gpc1_1 gpc1_1_668(
      {stage064[28]},
      {stage064[82]}
   );
   gpc1_1 gpc1_1_669(
      {stage064[29]},
      {stage064[83]}
   );
   gpc1_1 gpc1_1_670(
      {stage064[30]},
      {stage064[84]}
   );
   gpc1_1 gpc1_1_671(
      {stage064[31]},
      {stage064[85]}
   );
   gpc1_1 gpc1_1_672(
      {stage064[32]},
      {stage064[86]}
   );
   gpc1_1 gpc1_1_673(
      {stage064[33]},
      {stage064[87]}
   );
   gpc1_1 gpc1_1_674(
      {stage064[34]},
      {stage064[88]}
   );
   gpc1_1 gpc1_1_675(
      {stage064[35]},
      {stage064[89]}
   );
   gpc1_1 gpc1_1_676(
      {stage064[36]},
      {stage064[90]}
   );
   gpc1_1 gpc1_1_677(
      {stage064[37]},
      {stage064[91]}
   );
   gpc1_1 gpc1_1_678(
      {stage064[38]},
      {stage064[92]}
   );
   gpc606_5 gpc606_5_679(
      {stage064[39], stage064[40], stage064[41], stage064[42], stage064[43], stage064[44]},
      {stage066[0], stage066[1], stage066[2], stage066[3], stage066[4], stage066[5]},
      {stage068[59], stage067[67], stage066[72], stage065[73], stage064[93]}
   );
   gpc606_5 gpc606_5_680(
      {stage064[45], stage064[46], stage064[47], stage064[48], stage064[49], stage064[50]},
      {stage066[6], stage066[7], stage066[8], stage066[9], stage066[10], stage066[11]},
      {stage068[60], stage067[68], stage066[73], stage065[74], stage064[94]}
   );
   gpc606_5 gpc606_5_681(
      {stage064[51], stage064[52], stage064[53], stage064[54], stage064[55], stage064[56]},
      {stage066[12], stage066[13], stage066[14], stage066[15], stage066[16], stage066[17]},
      {stage068[61], stage067[69], stage066[74], stage065[75], stage064[95]}
   );
   gpc606_5 gpc606_5_682(
      {stage064[57], stage064[58], stage064[59], stage064[60], stage064[61], stage064[62]},
      {stage066[18], stage066[19], stage066[20], stage066[21], stage066[22], stage066[23]},
      {stage068[62], stage067[70], stage066[75], stage065[76], stage064[96]}
   );
   gpc1_1 gpc1_1_683(
      {stage065[42]},
      {stage065[77]}
   );
   gpc1_1 gpc1_1_684(
      {stage065[43]},
      {stage065[78]}
   );
   gpc1_1 gpc1_1_685(
      {stage065[44]},
      {stage065[79]}
   );
   gpc1_1 gpc1_1_686(
      {stage065[45]},
      {stage065[80]}
   );
   gpc1_1 gpc1_1_687(
      {stage065[46]},
      {stage065[81]}
   );
   gpc1_1 gpc1_1_688(
      {stage065[47]},
      {stage065[82]}
   );
   gpc1_1 gpc1_1_689(
      {stage065[48]},
      {stage065[83]}
   );
   gpc1_1 gpc1_1_690(
      {stage065[49]},
      {stage065[84]}
   );
   gpc1_1 gpc1_1_691(
      {stage065[50]},
      {stage065[85]}
   );
   gpc1_1 gpc1_1_692(
      {stage065[51]},
      {stage065[86]}
   );
   gpc1_1 gpc1_1_693(
      {stage065[52]},
      {stage065[87]}
   );
   gpc623_5 gpc623_5_694(
      {stage065[53], stage065[54], stage065[55]},
      {stage066[24], stage066[25]},
      {stage067[0], stage067[1], stage067[2], stage067[3], stage067[4], stage067[5]},
      {stage069[58], stage068[63], stage067[71], stage066[76], stage065[88]}
   );
   gpc623_5 gpc623_5_695(
      {stage065[56], stage065[57], stage065[58]},
      {stage066[26], stage066[27]},
      {stage067[6], stage067[7], stage067[8], stage067[9], stage067[10], stage067[11]},
      {stage069[59], stage068[64], stage067[72], stage066[77], stage065[89]}
   );
   gpc623_5 gpc623_5_696(
      {stage065[59], stage065[60], stage065[61]},
      {stage066[28], stage066[29]},
      {stage067[12], stage067[13], stage067[14], stage067[15], stage067[16], stage067[17]},
      {stage069[60], stage068[65], stage067[73], stage066[78], stage065[90]}
   );
   gpc1_1 gpc1_1_697(
      {stage066[30]},
      {stage066[79]}
   );
   gpc606_5 gpc606_5_698(
      {stage066[31], stage066[32], stage066[33], stage066[34], stage066[35], stage066[36]},
      {stage068[0], stage068[1], stage068[2], stage068[3], stage068[4], stage068[5]},
      {stage070[57], stage069[61], stage068[66], stage067[74], stage066[80]}
   );
   gpc606_5 gpc606_5_699(
      {stage066[37], stage066[38], stage066[39], stage066[40], stage066[41], stage066[42]},
      {stage068[6], stage068[7], stage068[8], stage068[9], stage068[10], stage068[11]},
      {stage070[58], stage069[62], stage068[67], stage067[75], stage066[81]}
   );
   gpc606_5 gpc606_5_700(
      {stage066[43], stage066[44], stage066[45], stage066[46], stage066[47], stage066[48]},
      {stage068[12], stage068[13], stage068[14], stage068[15], stage068[16], stage068[17]},
      {stage070[59], stage069[63], stage068[68], stage067[76], stage066[82]}
   );
   gpc606_5 gpc606_5_701(
      {stage066[49], stage066[50], stage066[51], stage066[52], stage066[53], stage066[54]},
      {stage068[18], stage068[19], stage068[20], stage068[21], stage068[22], stage068[23]},
      {stage070[60], stage069[64], stage068[69], stage067[77], stage066[83]}
   );
   gpc606_5 gpc606_5_702(
      {stage066[55], stage066[56], stage066[57], stage066[58], stage066[59], stage066[60]},
      {stage068[24], stage068[25], stage068[26], stage068[27], stage068[28], stage068[29]},
      {stage070[61], stage069[65], stage068[70], stage067[78], stage066[84]}
   );
   gpc1_1 gpc1_1_703(
      {stage067[18]},
      {stage067[79]}
   );
   gpc1_1 gpc1_1_704(
      {stage067[19]},
      {stage067[80]}
   );
   gpc1_1 gpc1_1_705(
      {stage067[20]},
      {stage067[81]}
   );
   gpc1_1 gpc1_1_706(
      {stage067[21]},
      {stage067[82]}
   );
   gpc1_1 gpc1_1_707(
      {stage067[22]},
      {stage067[83]}
   );
   gpc1_1 gpc1_1_708(
      {stage067[23]},
      {stage067[84]}
   );
   gpc1_1 gpc1_1_709(
      {stage067[24]},
      {stage067[85]}
   );
   gpc1_1 gpc1_1_710(
      {stage067[25]},
      {stage067[86]}
   );
   gpc1_1 gpc1_1_711(
      {stage067[26]},
      {stage067[87]}
   );
   gpc1_1 gpc1_1_712(
      {stage067[27]},
      {stage067[88]}
   );
   gpc1_1 gpc1_1_713(
      {stage067[28]},
      {stage067[89]}
   );
   gpc1_1 gpc1_1_714(
      {stage067[29]},
      {stage067[90]}
   );
   gpc1_1 gpc1_1_715(
      {stage067[30]},
      {stage067[91]}
   );
   gpc1_1 gpc1_1_716(
      {stage067[31]},
      {stage067[92]}
   );
   gpc1_1 gpc1_1_717(
      {stage067[32]},
      {stage067[93]}
   );
   gpc1_1 gpc1_1_718(
      {stage067[33]},
      {stage067[94]}
   );
   gpc1_1 gpc1_1_719(
      {stage067[34]},
      {stage067[95]}
   );
   gpc1_1 gpc1_1_720(
      {stage067[35]},
      {stage067[96]}
   );
   gpc1_1 gpc1_1_721(
      {stage067[36]},
      {stage067[97]}
   );
   gpc1_1 gpc1_1_722(
      {stage067[37]},
      {stage067[98]}
   );
   gpc615_5 gpc615_5_723(
      {stage067[38], stage067[39], stage067[40], stage067[41], stage067[42]},
      {stage068[30]},
      {stage069[0], stage069[1], stage069[2], stage069[3], stage069[4], stage069[5]},
      {stage071[56], stage070[62], stage069[66], stage068[71], stage067[99]}
   );
   gpc615_5 gpc615_5_724(
      {stage067[43], stage067[44], stage067[45], stage067[46], stage067[47]},
      {stage068[31]},
      {stage069[6], stage069[7], stage069[8], stage069[9], stage069[10], stage069[11]},
      {stage071[57], stage070[63], stage069[67], stage068[72], stage067[100]}
   );
   gpc615_5 gpc615_5_725(
      {stage067[48], stage067[49], stage067[50], stage067[51], stage067[52]},
      {stage068[32]},
      {stage069[12], stage069[13], stage069[14], stage069[15], stage069[16], stage069[17]},
      {stage071[58], stage070[64], stage069[68], stage068[73], stage067[101]}
   );
   gpc207_4 gpc207_4_726(
      {stage067[53], stage067[54], stage067[55], stage067[56], stage067[57], stage067[58], stage067[59]},
      {stage069[18], stage069[19]},
      {stage070[65], stage069[69], stage068[74], stage067[102]}
   );
   gpc1_1 gpc1_1_727(
      {stage068[33]},
      {stage068[75]}
   );
   gpc1_1 gpc1_1_728(
      {stage068[34]},
      {stage068[76]}
   );
   gpc1_1 gpc1_1_729(
      {stage068[35]},
      {stage068[77]}
   );
   gpc1_1 gpc1_1_730(
      {stage068[36]},
      {stage068[78]}
   );
   gpc1_1 gpc1_1_731(
      {stage068[37]},
      {stage068[79]}
   );
   gpc1_1 gpc1_1_732(
      {stage068[38]},
      {stage068[80]}
   );
   gpc615_5 gpc615_5_733(
      {stage068[39], stage068[40], stage068[41], stage068[42], stage068[43]},
      {stage069[20]},
      {stage070[0], stage070[1], stage070[2], stage070[3], stage070[4], stage070[5]},
      {stage072[55], stage071[59], stage070[66], stage069[70], stage068[81]}
   );
   gpc615_5 gpc615_5_734(
      {stage068[44], stage068[45], stage068[46], stage068[47], stage068[48]},
      {stage069[21]},
      {stage070[6], stage070[7], stage070[8], stage070[9], stage070[10], stage070[11]},
      {stage072[56], stage071[60], stage070[67], stage069[71], stage068[82]}
   );
   gpc615_5 gpc615_5_735(
      {stage068[49], stage068[50], stage068[51], stage068[52], stage068[53]},
      {stage069[22]},
      {stage070[12], stage070[13], stage070[14], stage070[15], stage070[16], stage070[17]},
      {stage072[57], stage071[61], stage070[68], stage069[72], stage068[83]}
   );
   gpc615_5 gpc615_5_736(
      {stage068[54], stage068[55], stage068[56], stage068[57], stage068[58]},
      {stage069[23]},
      {stage070[18], stage070[19], stage070[20], stage070[21], stage070[22], stage070[23]},
      {stage072[58], stage071[62], stage070[69], stage069[73], stage068[84]}
   );
   gpc1_1 gpc1_1_737(
      {stage069[24]},
      {stage069[74]}
   );
   gpc1_1 gpc1_1_738(
      {stage069[25]},
      {stage069[75]}
   );
   gpc1_1 gpc1_1_739(
      {stage069[26]},
      {stage069[76]}
   );
   gpc1_1 gpc1_1_740(
      {stage069[27]},
      {stage069[77]}
   );
   gpc1_1 gpc1_1_741(
      {stage069[28]},
      {stage069[78]}
   );
   gpc1_1 gpc1_1_742(
      {stage069[29]},
      {stage069[79]}
   );
   gpc1_1 gpc1_1_743(
      {stage069[30]},
      {stage069[80]}
   );
   gpc1_1 gpc1_1_744(
      {stage069[31]},
      {stage069[81]}
   );
   gpc1_1 gpc1_1_745(
      {stage069[32]},
      {stage069[82]}
   );
   gpc1_1 gpc1_1_746(
      {stage069[33]},
      {stage069[83]}
   );
   gpc1_1 gpc1_1_747(
      {stage069[34]},
      {stage069[84]}
   );
   gpc1_1 gpc1_1_748(
      {stage069[35]},
      {stage069[85]}
   );
   gpc1_1 gpc1_1_749(
      {stage069[36]},
      {stage069[86]}
   );
   gpc1_1 gpc1_1_750(
      {stage069[37]},
      {stage069[87]}
   );
   gpc615_5 gpc615_5_751(
      {stage069[38], stage069[39], stage069[40], stage069[41], stage069[42]},
      {stage070[24]},
      {stage071[0], stage071[1], stage071[2], stage071[3], stage071[4], stage071[5]},
      {stage073[54], stage072[59], stage071[63], stage070[70], stage069[88]}
   );
   gpc615_5 gpc615_5_752(
      {stage069[43], stage069[44], stage069[45], stage069[46], stage069[47]},
      {stage070[25]},
      {stage071[6], stage071[7], stage071[8], stage071[9], stage071[10], stage071[11]},
      {stage073[55], stage072[60], stage071[64], stage070[71], stage069[89]}
   );
   gpc615_5 gpc615_5_753(
      {stage069[48], stage069[49], stage069[50], stage069[51], stage069[52]},
      {stage070[26]},
      {stage071[12], stage071[13], stage071[14], stage071[15], stage071[16], stage071[17]},
      {stage073[56], stage072[61], stage071[65], stage070[72], stage069[90]}
   );
   gpc615_5 gpc615_5_754(
      {stage069[53], stage069[54], stage069[55], stage069[56], stage069[57]},
      {stage070[27]},
      {stage071[18], stage071[19], stage071[20], stage071[21], stage071[22], stage071[23]},
      {stage073[57], stage072[62], stage071[66], stage070[73], stage069[91]}
   );
   gpc1_1 gpc1_1_755(
      {stage070[28]},
      {stage070[74]}
   );
   gpc1_1 gpc1_1_756(
      {stage070[29]},
      {stage070[75]}
   );
   gpc1_1 gpc1_1_757(
      {stage070[30]},
      {stage070[76]}
   );
   gpc1_1 gpc1_1_758(
      {stage070[31]},
      {stage070[77]}
   );
   gpc1_1 gpc1_1_759(
      {stage070[32]},
      {stage070[78]}
   );
   gpc1_1 gpc1_1_760(
      {stage070[33]},
      {stage070[79]}
   );
   gpc1_1 gpc1_1_761(
      {stage070[34]},
      {stage070[80]}
   );
   gpc1_1 gpc1_1_762(
      {stage070[35]},
      {stage070[81]}
   );
   gpc1_1 gpc1_1_763(
      {stage070[36]},
      {stage070[82]}
   );
   gpc1_1 gpc1_1_764(
      {stage070[37]},
      {stage070[83]}
   );
   gpc1_1 gpc1_1_765(
      {stage070[38]},
      {stage070[84]}
   );
   gpc1_1 gpc1_1_766(
      {stage070[39]},
      {stage070[85]}
   );
   gpc1_1 gpc1_1_767(
      {stage070[40]},
      {stage070[86]}
   );
   gpc606_5 gpc606_5_768(
      {stage070[41], stage070[42], stage070[43], stage070[44], stage070[45], stage070[46]},
      {stage072[0], stage072[1], stage072[2], stage072[3], stage072[4], stage072[5]},
      {stage074[53], stage073[58], stage072[63], stage071[67], stage070[87]}
   );
   gpc615_5 gpc615_5_769(
      {stage070[47], stage070[48], stage070[49], stage070[50], stage070[51]},
      {stage071[24]},
      {stage072[6], stage072[7], stage072[8], stage072[9], stage072[10], stage072[11]},
      {stage074[54], stage073[59], stage072[64], stage071[68], stage070[88]}
   );
   gpc615_5 gpc615_5_770(
      {stage070[52], stage070[53], stage070[54], stage070[55], stage070[56]},
      {stage071[25]},
      {stage072[12], stage072[13], stage072[14], stage072[15], stage072[16], stage072[17]},
      {stage074[55], stage073[60], stage072[65], stage071[69], stage070[89]}
   );
   gpc1_1 gpc1_1_771(
      {stage071[26]},
      {stage071[70]}
   );
   gpc1_1 gpc1_1_772(
      {stage071[27]},
      {stage071[71]}
   );
   gpc1_1 gpc1_1_773(
      {stage071[28]},
      {stage071[72]}
   );
   gpc1_1 gpc1_1_774(
      {stage071[29]},
      {stage071[73]}
   );
   gpc1_1 gpc1_1_775(
      {stage071[30]},
      {stage071[74]}
   );
   gpc615_5 gpc615_5_776(
      {stage071[31], stage071[32], stage071[33], stage071[34], stage071[35]},
      {stage072[18]},
      {stage073[0], stage073[1], stage073[2], stage073[3], stage073[4], stage073[5]},
      {stage075[52], stage074[56], stage073[61], stage072[66], stage071[75]}
   );
   gpc615_5 gpc615_5_777(
      {stage071[36], stage071[37], stage071[38], stage071[39], stage071[40]},
      {stage072[19]},
      {stage073[6], stage073[7], stage073[8], stage073[9], stage073[10], stage073[11]},
      {stage075[53], stage074[57], stage073[62], stage072[67], stage071[76]}
   );
   gpc615_5 gpc615_5_778(
      {stage071[41], stage071[42], stage071[43], stage071[44], stage071[45]},
      {stage072[20]},
      {stage073[12], stage073[13], stage073[14], stage073[15], stage073[16], stage073[17]},
      {stage075[54], stage074[58], stage073[63], stage072[68], stage071[77]}
   );
   gpc615_5 gpc615_5_779(
      {stage071[46], stage071[47], stage071[48], stage071[49], stage071[50]},
      {stage072[21]},
      {stage073[18], stage073[19], stage073[20], stage073[21], stage073[22], stage073[23]},
      {stage075[55], stage074[59], stage073[64], stage072[69], stage071[78]}
   );
   gpc615_5 gpc615_5_780(
      {stage071[51], stage071[52], stage071[53], stage071[54], stage071[55]},
      {stage072[22]},
      {stage073[24], stage073[25], stage073[26], stage073[27], stage073[28], stage073[29]},
      {stage075[56], stage074[60], stage073[65], stage072[70], stage071[79]}
   );
   gpc1_1 gpc1_1_781(
      {stage072[23]},
      {stage072[71]}
   );
   gpc1_1 gpc1_1_782(
      {stage072[24]},
      {stage072[72]}
   );
   gpc1_1 gpc1_1_783(
      {stage072[25]},
      {stage072[73]}
   );
   gpc1_1 gpc1_1_784(
      {stage072[26]},
      {stage072[74]}
   );
   gpc1_1 gpc1_1_785(
      {stage072[27]},
      {stage072[75]}
   );
   gpc1_1 gpc1_1_786(
      {stage072[28]},
      {stage072[76]}
   );
   gpc1_1 gpc1_1_787(
      {stage072[29]},
      {stage072[77]}
   );
   gpc1_1 gpc1_1_788(
      {stage072[30]},
      {stage072[78]}
   );
   gpc606_5 gpc606_5_789(
      {stage072[31], stage072[32], stage072[33], stage072[34], stage072[35], stage072[36]},
      {stage074[0], stage074[1], stage074[2], stage074[3], stage074[4], stage074[5]},
      {stage076[51], stage075[57], stage074[61], stage073[66], stage072[79]}
   );
   gpc606_5 gpc606_5_790(
      {stage072[37], stage072[38], stage072[39], stage072[40], stage072[41], stage072[42]},
      {stage074[6], stage074[7], stage074[8], stage074[9], stage074[10], stage074[11]},
      {stage076[52], stage075[58], stage074[62], stage073[67], stage072[80]}
   );
   gpc606_5 gpc606_5_791(
      {stage072[43], stage072[44], stage072[45], stage072[46], stage072[47], stage072[48]},
      {stage074[12], stage074[13], stage074[14], stage074[15], stage074[16], stage074[17]},
      {stage076[53], stage075[59], stage074[63], stage073[68], stage072[81]}
   );
   gpc606_5 gpc606_5_792(
      {stage072[49], stage072[50], stage072[51], stage072[52], stage072[53], stage072[54]},
      {stage074[18], stage074[19], stage074[20], stage074[21], stage074[22], stage074[23]},
      {stage076[54], stage075[60], stage074[64], stage073[69], stage072[82]}
   );
   gpc1_1 gpc1_1_793(
      {stage073[30]},
      {stage073[70]}
   );
   gpc1_1 gpc1_1_794(
      {stage073[31]},
      {stage073[71]}
   );
   gpc1_1 gpc1_1_795(
      {stage073[32]},
      {stage073[72]}
   );
   gpc1_1 gpc1_1_796(
      {stage073[33]},
      {stage073[73]}
   );
   gpc1_1 gpc1_1_797(
      {stage073[34]},
      {stage073[74]}
   );
   gpc1_1 gpc1_1_798(
      {stage073[35]},
      {stage073[75]}
   );
   gpc1_1 gpc1_1_799(
      {stage073[36]},
      {stage073[76]}
   );
   gpc1_1 gpc1_1_800(
      {stage073[37]},
      {stage073[77]}
   );
   gpc1_1 gpc1_1_801(
      {stage073[38]},
      {stage073[78]}
   );
   gpc1_1 gpc1_1_802(
      {stage073[39]},
      {stage073[79]}
   );
   gpc1_1 gpc1_1_803(
      {stage073[40]},
      {stage073[80]}
   );
   gpc1_1 gpc1_1_804(
      {stage073[41]},
      {stage073[81]}
   );
   gpc606_5 gpc606_5_805(
      {stage073[42], stage073[43], stage073[44], stage073[45], stage073[46], stage073[47]},
      {stage075[0], stage075[1], stage075[2], stage075[3], stage075[4], stage075[5]},
      {stage077[50], stage076[55], stage075[61], stage074[65], stage073[82]}
   );
   gpc606_5 gpc606_5_806(
      {stage073[48], stage073[49], stage073[50], stage073[51], stage073[52], stage073[53]},
      {stage075[6], stage075[7], stage075[8], stage075[9], stage075[10], stage075[11]},
      {stage077[51], stage076[56], stage075[62], stage074[66], stage073[83]}
   );
   gpc1_1 gpc1_1_807(
      {stage074[24]},
      {stage074[67]}
   );
   gpc1_1 gpc1_1_808(
      {stage074[25]},
      {stage074[68]}
   );
   gpc1_1 gpc1_1_809(
      {stage074[26]},
      {stage074[69]}
   );
   gpc1_1 gpc1_1_810(
      {stage074[27]},
      {stage074[70]}
   );
   gpc1_1 gpc1_1_811(
      {stage074[28]},
      {stage074[71]}
   );
   gpc1_1 gpc1_1_812(
      {stage074[29]},
      {stage074[72]}
   );
   gpc1_1 gpc1_1_813(
      {stage074[30]},
      {stage074[73]}
   );
   gpc1_1 gpc1_1_814(
      {stage074[31]},
      {stage074[74]}
   );
   gpc1_1 gpc1_1_815(
      {stage074[32]},
      {stage074[75]}
   );
   gpc1_1 gpc1_1_816(
      {stage074[33]},
      {stage074[76]}
   );
   gpc1_1 gpc1_1_817(
      {stage074[34]},
      {stage074[77]}
   );
   gpc606_5 gpc606_5_818(
      {stage074[35], stage074[36], stage074[37], stage074[38], stage074[39], stage074[40]},
      {stage076[0], stage076[1], stage076[2], stage076[3], stage076[4], stage076[5]},
      {stage078[49], stage077[52], stage076[57], stage075[63], stage074[78]}
   );
   gpc606_5 gpc606_5_819(
      {stage074[41], stage074[42], stage074[43], stage074[44], stage074[45], stage074[46]},
      {stage076[6], stage076[7], stage076[8], stage076[9], stage076[10], stage076[11]},
      {stage078[50], stage077[53], stage076[58], stage075[64], stage074[79]}
   );
   gpc606_5 gpc606_5_820(
      {stage074[47], stage074[48], stage074[49], stage074[50], stage074[51], stage074[52]},
      {stage076[12], stage076[13], stage076[14], stage076[15], stage076[16], stage076[17]},
      {stage078[51], stage077[54], stage076[59], stage075[65], stage074[80]}
   );
   gpc1_1 gpc1_1_821(
      {stage075[12]},
      {stage075[66]}
   );
   gpc1_1 gpc1_1_822(
      {stage075[13]},
      {stage075[67]}
   );
   gpc1_1 gpc1_1_823(
      {stage075[14]},
      {stage075[68]}
   );
   gpc1_1 gpc1_1_824(
      {stage075[15]},
      {stage075[69]}
   );
   gpc1_1 gpc1_1_825(
      {stage075[16]},
      {stage075[70]}
   );
   gpc1_1 gpc1_1_826(
      {stage075[17]},
      {stage075[71]}
   );
   gpc606_5 gpc606_5_827(
      {stage075[18], stage075[19], stage075[20], stage075[21], stage075[22], stage075[23]},
      {stage077[0], stage077[1], stage077[2], stage077[3], stage077[4], stage077[5]},
      {stage079[48], stage078[52], stage077[55], stage076[60], stage075[72]}
   );
   gpc606_5 gpc606_5_828(
      {stage075[24], stage075[25], stage075[26], stage075[27], stage075[28], stage075[29]},
      {stage077[6], stage077[7], stage077[8], stage077[9], stage077[10], stage077[11]},
      {stage079[49], stage078[53], stage077[56], stage076[61], stage075[73]}
   );
   gpc606_5 gpc606_5_829(
      {stage075[30], stage075[31], stage075[32], stage075[33], stage075[34], stage075[35]},
      {stage077[12], stage077[13], stage077[14], stage077[15], stage077[16], stage077[17]},
      {stage079[50], stage078[54], stage077[57], stage076[62], stage075[74]}
   );
   gpc606_5 gpc606_5_830(
      {stage075[36], stage075[37], stage075[38], stage075[39], stage075[40], stage075[41]},
      {stage077[18], stage077[19], stage077[20], stage077[21], stage077[22], stage077[23]},
      {stage079[51], stage078[55], stage077[58], stage076[63], stage075[75]}
   );
   gpc2135_5 gpc2135_5_831(
      {stage075[42], stage075[43], stage075[44], stage075[45], stage075[46]},
      {stage076[18], stage076[19], stage076[20]},
      {stage077[24]},
      {stage078[0], stage078[1]},
      {stage079[52], stage078[56], stage077[59], stage076[64], stage075[76]}
   );
   gpc2135_5 gpc2135_5_832(
      {stage075[47], stage075[48], stage075[49], stage075[50], stage075[51]},
      {stage076[21], stage076[22], stage076[23]},
      {stage077[25]},
      {stage078[2], stage078[3]},
      {stage079[53], stage078[57], stage077[60], stage076[65], stage075[77]}
   );
   gpc1_1 gpc1_1_833(
      {stage076[24]},
      {stage076[66]}
   );
   gpc1_1 gpc1_1_834(
      {stage076[25]},
      {stage076[67]}
   );
   gpc1_1 gpc1_1_835(
      {stage076[26]},
      {stage076[68]}
   );
   gpc606_5 gpc606_5_836(
      {stage076[27], stage076[28], stage076[29], stage076[30], stage076[31], stage076[32]},
      {stage078[4], stage078[5], stage078[6], stage078[7], stage078[8], stage078[9]},
      {stage080[47], stage079[54], stage078[58], stage077[61], stage076[69]}
   );
   gpc606_5 gpc606_5_837(
      {stage076[33], stage076[34], stage076[35], stage076[36], stage076[37], stage076[38]},
      {stage078[10], stage078[11], stage078[12], stage078[13], stage078[14], stage078[15]},
      {stage080[48], stage079[55], stage078[59], stage077[62], stage076[70]}
   );
   gpc606_5 gpc606_5_838(
      {stage076[39], stage076[40], stage076[41], stage076[42], stage076[43], stage076[44]},
      {stage078[16], stage078[17], stage078[18], stage078[19], stage078[20], stage078[21]},
      {stage080[49], stage079[56], stage078[60], stage077[63], stage076[71]}
   );
   gpc606_5 gpc606_5_839(
      {stage076[45], stage076[46], stage076[47], stage076[48], stage076[49], stage076[50]},
      {stage078[22], stage078[23], stage078[24], stage078[25], stage078[26], stage078[27]},
      {stage080[50], stage079[57], stage078[61], stage077[64], stage076[72]}
   );
   gpc1_1 gpc1_1_840(
      {stage077[26]},
      {stage077[65]}
   );
   gpc1_1 gpc1_1_841(
      {stage077[27]},
      {stage077[66]}
   );
   gpc1_1 gpc1_1_842(
      {stage077[28]},
      {stage077[67]}
   );
   gpc1_1 gpc1_1_843(
      {stage077[29]},
      {stage077[68]}
   );
   gpc1_1 gpc1_1_844(
      {stage077[30]},
      {stage077[69]}
   );
   gpc1_1 gpc1_1_845(
      {stage077[31]},
      {stage077[70]}
   );
   gpc1_1 gpc1_1_846(
      {stage077[32]},
      {stage077[71]}
   );
   gpc606_5 gpc606_5_847(
      {stage077[33], stage077[34], stage077[35], stage077[36], stage077[37], stage077[38]},
      {stage079[0], stage079[1], stage079[2], stage079[3], stage079[4], stage079[5]},
      {stage081[46], stage080[51], stage079[58], stage078[62], stage077[72]}
   );
   gpc606_5 gpc606_5_848(
      {stage077[39], stage077[40], stage077[41], stage077[42], stage077[43], stage077[44]},
      {stage079[6], stage079[7], stage079[8], stage079[9], stage079[10], stage079[11]},
      {stage081[47], stage080[52], stage079[59], stage078[63], stage077[73]}
   );
   gpc615_5 gpc615_5_849(
      {stage077[45], stage077[46], stage077[47], stage077[48], stage077[49]},
      {stage078[28]},
      {stage079[12], stage079[13], stage079[14], stage079[15], stage079[16], stage079[17]},
      {stage081[48], stage080[53], stage079[60], stage078[64], stage077[74]}
   );
   gpc1_1 gpc1_1_850(
      {stage078[29]},
      {stage078[65]}
   );
   gpc1_1 gpc1_1_851(
      {stage078[30]},
      {stage078[66]}
   );
   gpc1_1 gpc1_1_852(
      {stage078[31]},
      {stage078[67]}
   );
   gpc606_5 gpc606_5_853(
      {stage078[32], stage078[33], stage078[34], stage078[35], stage078[36], stage078[37]},
      {stage080[0], stage080[1], stage080[2], stage080[3], stage080[4], stage080[5]},
      {stage082[45], stage081[49], stage080[54], stage079[61], stage078[68]}
   );
   gpc606_5 gpc606_5_854(
      {stage078[38], stage078[39], stage078[40], stage078[41], stage078[42], stage078[43]},
      {stage080[6], stage080[7], stage080[8], stage080[9], stage080[10], stage080[11]},
      {stage082[46], stage081[50], stage080[55], stage079[62], stage078[69]}
   );
   gpc615_5 gpc615_5_855(
      {stage078[44], stage078[45], stage078[46], stage078[47], stage078[48]},
      {stage079[18]},
      {stage080[12], stage080[13], stage080[14], stage080[15], stage080[16], stage080[17]},
      {stage082[47], stage081[51], stage080[56], stage079[63], stage078[70]}
   );
   gpc1_1 gpc1_1_856(
      {stage079[19]},
      {stage079[64]}
   );
   gpc1_1 gpc1_1_857(
      {stage079[20]},
      {stage079[65]}
   );
   gpc1_1 gpc1_1_858(
      {stage079[21]},
      {stage079[66]}
   );
   gpc1_1 gpc1_1_859(
      {stage079[22]},
      {stage079[67]}
   );
   gpc1_1 gpc1_1_860(
      {stage079[23]},
      {stage079[68]}
   );
   gpc1_1 gpc1_1_861(
      {stage079[24]},
      {stage079[69]}
   );
   gpc1_1 gpc1_1_862(
      {stage079[25]},
      {stage079[70]}
   );
   gpc1_1 gpc1_1_863(
      {stage079[26]},
      {stage079[71]}
   );
   gpc1_1 gpc1_1_864(
      {stage079[27]},
      {stage079[72]}
   );
   gpc1_1 gpc1_1_865(
      {stage079[28]},
      {stage079[73]}
   );
   gpc1_1 gpc1_1_866(
      {stage079[29]},
      {stage079[74]}
   );
   gpc1_1 gpc1_1_867(
      {stage079[30]},
      {stage079[75]}
   );
   gpc1_1 gpc1_1_868(
      {stage079[31]},
      {stage079[76]}
   );
   gpc1_1 gpc1_1_869(
      {stage079[32]},
      {stage079[77]}
   );
   gpc1_1 gpc1_1_870(
      {stage079[33]},
      {stage079[78]}
   );
   gpc1_1 gpc1_1_871(
      {stage079[34]},
      {stage079[79]}
   );
   gpc1_1 gpc1_1_872(
      {stage079[35]},
      {stage079[80]}
   );
   gpc1_1 gpc1_1_873(
      {stage079[36]},
      {stage079[81]}
   );
   gpc1_1 gpc1_1_874(
      {stage079[37]},
      {stage079[82]}
   );
   gpc615_5 gpc615_5_875(
      {stage079[38], stage079[39], stage079[40], stage079[41], stage079[42]},
      {stage080[18]},
      {stage081[0], stage081[1], stage081[2], stage081[3], stage081[4], stage081[5]},
      {stage083[44], stage082[48], stage081[52], stage080[57], stage079[83]}
   );
   gpc615_5 gpc615_5_876(
      {stage079[43], stage079[44], stage079[45], stage079[46], stage079[47]},
      {stage080[19]},
      {stage081[6], stage081[7], stage081[8], stage081[9], stage081[10], stage081[11]},
      {stage083[45], stage082[49], stage081[53], stage080[58], stage079[84]}
   );
   gpc1_1 gpc1_1_877(
      {stage080[20]},
      {stage080[59]}
   );
   gpc1_1 gpc1_1_878(
      {stage080[21]},
      {stage080[60]}
   );
   gpc1_1 gpc1_1_879(
      {stage080[22]},
      {stage080[61]}
   );
   gpc1_1 gpc1_1_880(
      {stage080[23]},
      {stage080[62]}
   );
   gpc1_1 gpc1_1_881(
      {stage080[24]},
      {stage080[63]}
   );
   gpc1_1 gpc1_1_882(
      {stage080[25]},
      {stage080[64]}
   );
   gpc1_1 gpc1_1_883(
      {stage080[26]},
      {stage080[65]}
   );
   gpc1_1 gpc1_1_884(
      {stage080[27]},
      {stage080[66]}
   );
   gpc1_1 gpc1_1_885(
      {stage080[28]},
      {stage080[67]}
   );
   gpc606_5 gpc606_5_886(
      {stage080[29], stage080[30], stage080[31], stage080[32], stage080[33], stage080[34]},
      {stage082[0], stage082[1], stage082[2], stage082[3], stage082[4], stage082[5]},
      {stage084[43], stage083[46], stage082[50], stage081[54], stage080[68]}
   );
   gpc606_5 gpc606_5_887(
      {stage080[35], stage080[36], stage080[37], stage080[38], stage080[39], stage080[40]},
      {stage082[6], stage082[7], stage082[8], stage082[9], stage082[10], stage082[11]},
      {stage084[44], stage083[47], stage082[51], stage081[55], stage080[69]}
   );
   gpc606_5 gpc606_5_888(
      {stage080[41], stage080[42], stage080[43], stage080[44], stage080[45], stage080[46]},
      {stage082[12], stage082[13], stage082[14], stage082[15], stage082[16], stage082[17]},
      {stage084[45], stage083[48], stage082[52], stage081[56], stage080[70]}
   );
   gpc1_1 gpc1_1_889(
      {stage081[12]},
      {stage081[57]}
   );
   gpc1_1 gpc1_1_890(
      {stage081[13]},
      {stage081[58]}
   );
   gpc1_1 gpc1_1_891(
      {stage081[14]},
      {stage081[59]}
   );
   gpc1_1 gpc1_1_892(
      {stage081[15]},
      {stage081[60]}
   );
   gpc1_1 gpc1_1_893(
      {stage081[16]},
      {stage081[61]}
   );
   gpc1_1 gpc1_1_894(
      {stage081[17]},
      {stage081[62]}
   );
   gpc1_1 gpc1_1_895(
      {stage081[18]},
      {stage081[63]}
   );
   gpc1_1 gpc1_1_896(
      {stage081[19]},
      {stage081[64]}
   );
   gpc1_1 gpc1_1_897(
      {stage081[20]},
      {stage081[65]}
   );
   gpc1_1 gpc1_1_898(
      {stage081[21]},
      {stage081[66]}
   );
   gpc1_1 gpc1_1_899(
      {stage081[22]},
      {stage081[67]}
   );
   gpc1_1 gpc1_1_900(
      {stage081[23]},
      {stage081[68]}
   );
   gpc1_1 gpc1_1_901(
      {stage081[24]},
      {stage081[69]}
   );
   gpc1_1 gpc1_1_902(
      {stage081[25]},
      {stage081[70]}
   );
   gpc615_5 gpc615_5_903(
      {stage081[26], stage081[27], stage081[28], stage081[29], stage081[30]},
      {stage082[18]},
      {stage083[0], stage083[1], stage083[2], stage083[3], stage083[4], stage083[5]},
      {stage085[42], stage084[46], stage083[49], stage082[53], stage081[71]}
   );
   gpc615_5 gpc615_5_904(
      {stage081[31], stage081[32], stage081[33], stage081[34], stage081[35]},
      {stage082[19]},
      {stage083[6], stage083[7], stage083[8], stage083[9], stage083[10], stage083[11]},
      {stage085[43], stage084[47], stage083[50], stage082[54], stage081[72]}
   );
   gpc615_5 gpc615_5_905(
      {stage081[36], stage081[37], stage081[38], stage081[39], stage081[40]},
      {stage082[20]},
      {stage083[12], stage083[13], stage083[14], stage083[15], stage083[16], stage083[17]},
      {stage085[44], stage084[48], stage083[51], stage082[55], stage081[73]}
   );
   gpc615_5 gpc615_5_906(
      {stage081[41], stage081[42], stage081[43], stage081[44], stage081[45]},
      {stage082[21]},
      {stage083[18], stage083[19], stage083[20], stage083[21], stage083[22], stage083[23]},
      {stage085[45], stage084[49], stage083[52], stage082[56], stage081[74]}
   );
   gpc1_1 gpc1_1_907(
      {stage082[22]},
      {stage082[57]}
   );
   gpc1_1 gpc1_1_908(
      {stage082[23]},
      {stage082[58]}
   );
   gpc1_1 gpc1_1_909(
      {stage082[24]},
      {stage082[59]}
   );
   gpc1_1 gpc1_1_910(
      {stage082[25]},
      {stage082[60]}
   );
   gpc1_1 gpc1_1_911(
      {stage082[26]},
      {stage082[61]}
   );
   gpc1_1 gpc1_1_912(
      {stage082[27]},
      {stage082[62]}
   );
   gpc606_5 gpc606_5_913(
      {stage082[28], stage082[29], stage082[30], stage082[31], stage082[32], stage082[33]},
      {stage084[0], stage084[1], stage084[2], stage084[3], stage084[4], stage084[5]},
      {stage086[41], stage085[46], stage084[50], stage083[53], stage082[63]}
   );
   gpc606_5 gpc606_5_914(
      {stage082[34], stage082[35], stage082[36], stage082[37], stage082[38], stage082[39]},
      {stage084[6], stage084[7], stage084[8], stage084[9], stage084[10], stage084[11]},
      {stage086[42], stage085[47], stage084[51], stage083[54], stage082[64]}
   );
   gpc615_5 gpc615_5_915(
      {stage082[40], stage082[41], stage082[42], stage082[43], stage082[44]},
      {stage083[24]},
      {stage084[12], stage084[13], stage084[14], stage084[15], stage084[16], stage084[17]},
      {stage086[43], stage085[48], stage084[52], stage083[55], stage082[65]}
   );
   gpc1_1 gpc1_1_916(
      {stage083[25]},
      {stage083[56]}
   );
   gpc1_1 gpc1_1_917(
      {stage083[26]},
      {stage083[57]}
   );
   gpc1_1 gpc1_1_918(
      {stage083[27]},
      {stage083[58]}
   );
   gpc1_1 gpc1_1_919(
      {stage083[28]},
      {stage083[59]}
   );
   gpc615_5 gpc615_5_920(
      {stage083[29], stage083[30], stage083[31], stage083[32], stage083[33]},
      {stage084[18]},
      {stage085[0], stage085[1], stage085[2], stage085[3], stage085[4], stage085[5]},
      {stage087[40], stage086[44], stage085[49], stage084[53], stage083[60]}
   );
   gpc615_5 gpc615_5_921(
      {stage083[34], stage083[35], stage083[36], stage083[37], stage083[38]},
      {stage084[19]},
      {stage085[6], stage085[7], stage085[8], stage085[9], stage085[10], stage085[11]},
      {stage087[41], stage086[45], stage085[50], stage084[54], stage083[61]}
   );
   gpc615_5 gpc615_5_922(
      {stage083[39], stage083[40], stage083[41], stage083[42], stage083[43]},
      {stage084[20]},
      {stage085[12], stage085[13], stage085[14], stage085[15], stage085[16], stage085[17]},
      {stage087[42], stage086[46], stage085[51], stage084[55], stage083[62]}
   );
   gpc1_1 gpc1_1_923(
      {stage084[21]},
      {stage084[56]}
   );
   gpc1_1 gpc1_1_924(
      {stage084[22]},
      {stage084[57]}
   );
   gpc1_1 gpc1_1_925(
      {stage084[23]},
      {stage084[58]}
   );
   gpc1_1 gpc1_1_926(
      {stage084[24]},
      {stage084[59]}
   );
   gpc1_1 gpc1_1_927(
      {stage084[25]},
      {stage084[60]}
   );
   gpc1_1 gpc1_1_928(
      {stage084[26]},
      {stage084[61]}
   );
   gpc1_1 gpc1_1_929(
      {stage084[27]},
      {stage084[62]}
   );
   gpc1_1 gpc1_1_930(
      {stage084[28]},
      {stage084[63]}
   );
   gpc1_1 gpc1_1_931(
      {stage084[29]},
      {stage084[64]}
   );
   gpc1_1 gpc1_1_932(
      {stage084[30]},
      {stage084[65]}
   );
   gpc1_1 gpc1_1_933(
      {stage084[31]},
      {stage084[66]}
   );
   gpc1_1 gpc1_1_934(
      {stage084[32]},
      {stage084[67]}
   );
   gpc1_1 gpc1_1_935(
      {stage084[33]},
      {stage084[68]}
   );
   gpc1_1 gpc1_1_936(
      {stage084[34]},
      {stage084[69]}
   );
   gpc1_1 gpc1_1_937(
      {stage084[35]},
      {stage084[70]}
   );
   gpc1_1 gpc1_1_938(
      {stage084[36]},
      {stage084[71]}
   );
   gpc1_1 gpc1_1_939(
      {stage084[37]},
      {stage084[72]}
   );
   gpc615_5 gpc615_5_940(
      {stage084[38], stage084[39], stage084[40], stage084[41], stage084[42]},
      {stage085[18]},
      {stage086[0], stage086[1], stage086[2], stage086[3], stage086[4], stage086[5]},
      {stage088[39], stage087[43], stage086[47], stage085[52], stage084[73]}
   );
   gpc1_1 gpc1_1_941(
      {stage085[19]},
      {stage085[53]}
   );
   gpc1_1 gpc1_1_942(
      {stage085[20]},
      {stage085[54]}
   );
   gpc1_1 gpc1_1_943(
      {stage085[21]},
      {stage085[55]}
   );
   gpc1_1 gpc1_1_944(
      {stage085[22]},
      {stage085[56]}
   );
   gpc1_1 gpc1_1_945(
      {stage085[23]},
      {stage085[57]}
   );
   gpc1_1 gpc1_1_946(
      {stage085[24]},
      {stage085[58]}
   );
   gpc1_1 gpc1_1_947(
      {stage085[25]},
      {stage085[59]}
   );
   gpc1_1 gpc1_1_948(
      {stage085[26]},
      {stage085[60]}
   );
   gpc1_1 gpc1_1_949(
      {stage085[27]},
      {stage085[61]}
   );
   gpc1_1 gpc1_1_950(
      {stage085[28]},
      {stage085[62]}
   );
   gpc1_1 gpc1_1_951(
      {stage085[29]},
      {stage085[63]}
   );
   gpc1_1 gpc1_1_952(
      {stage085[30]},
      {stage085[64]}
   );
   gpc1_1 gpc1_1_953(
      {stage085[31]},
      {stage085[65]}
   );
   gpc615_5 gpc615_5_954(
      {stage085[32], stage085[33], stage085[34], stage085[35], stage085[36]},
      {stage086[6]},
      {stage087[0], stage087[1], stage087[2], stage087[3], stage087[4], stage087[5]},
      {stage089[38], stage088[40], stage087[44], stage086[48], stage085[66]}
   );
   gpc615_5 gpc615_5_955(
      {stage085[37], stage085[38], stage085[39], stage085[40], stage085[41]},
      {stage086[7]},
      {stage087[6], stage087[7], stage087[8], stage087[9], stage087[10], stage087[11]},
      {stage089[39], stage088[41], stage087[45], stage086[49], stage085[67]}
   );
   gpc1_1 gpc1_1_956(
      {stage086[8]},
      {stage086[50]}
   );
   gpc1_1 gpc1_1_957(
      {stage086[9]},
      {stage086[51]}
   );
   gpc1_1 gpc1_1_958(
      {stage086[10]},
      {stage086[52]}
   );
   gpc1_1 gpc1_1_959(
      {stage086[11]},
      {stage086[53]}
   );
   gpc1_1 gpc1_1_960(
      {stage086[12]},
      {stage086[54]}
   );
   gpc1_1 gpc1_1_961(
      {stage086[13]},
      {stage086[55]}
   );
   gpc1_1 gpc1_1_962(
      {stage086[14]},
      {stage086[56]}
   );
   gpc1_1 gpc1_1_963(
      {stage086[15]},
      {stage086[57]}
   );
   gpc1_1 gpc1_1_964(
      {stage086[16]},
      {stage086[58]}
   );
   gpc1_1 gpc1_1_965(
      {stage086[17]},
      {stage086[59]}
   );
   gpc1_1 gpc1_1_966(
      {stage086[18]},
      {stage086[60]}
   );
   gpc1_1 gpc1_1_967(
      {stage086[19]},
      {stage086[61]}
   );
   gpc606_5 gpc606_5_968(
      {stage086[20], stage086[21], stage086[22], stage086[23], stage086[24], stage086[25]},
      {stage088[0], stage088[1], stage088[2], stage088[3], stage088[4], stage088[5]},
      {stage090[37], stage089[40], stage088[42], stage087[46], stage086[62]}
   );
   gpc606_5 gpc606_5_969(
      {stage086[26], stage086[27], stage086[28], stage086[29], stage086[30], stage086[31]},
      {stage088[6], stage088[7], stage088[8], stage088[9], stage088[10], stage088[11]},
      {stage090[38], stage089[41], stage088[43], stage087[47], stage086[63]}
   );
   gpc606_5 gpc606_5_970(
      {stage086[32], stage086[33], stage086[34], stage086[35], stage086[36], stage086[37]},
      {stage088[12], stage088[13], stage088[14], stage088[15], stage088[16], stage088[17]},
      {stage090[39], stage089[42], stage088[44], stage087[48], stage086[64]}
   );
   gpc1343_5 gpc1343_5_971(
      {stage086[38], stage086[39], stage086[40]},
      {stage087[12], stage087[13], stage087[14], stage087[15]},
      {stage088[18], stage088[19], stage088[20]},
      {stage089[0]},
      {stage090[40], stage089[43], stage088[45], stage087[49], stage086[65]}
   );
   gpc606_5 gpc606_5_972(
      {stage087[16], stage087[17], stage087[18], stage087[19], stage087[20], stage087[21]},
      {stage089[1], stage089[2], stage089[3], stage089[4], stage089[5], stage089[6]},
      {stage091[36], stage090[41], stage089[44], stage088[46], stage087[50]}
   );
   gpc606_5 gpc606_5_973(
      {stage087[22], stage087[23], stage087[24], stage087[25], stage087[26], stage087[27]},
      {stage089[7], stage089[8], stage089[9], stage089[10], stage089[11], stage089[12]},
      {stage091[37], stage090[42], stage089[45], stage088[47], stage087[51]}
   );
   gpc606_5 gpc606_5_974(
      {stage087[28], stage087[29], stage087[30], stage087[31], stage087[32], stage087[33]},
      {stage089[13], stage089[14], stage089[15], stage089[16], stage089[17], stage089[18]},
      {stage091[38], stage090[43], stage089[46], stage088[48], stage087[52]}
   );
   gpc606_5 gpc606_5_975(
      {stage087[34], stage087[35], stage087[36], stage087[37], stage087[38], stage087[39]},
      {stage089[19], stage089[20], stage089[21], stage089[22], stage089[23], stage089[24]},
      {stage091[39], stage090[44], stage089[47], stage088[49], stage087[53]}
   );
   gpc606_5 gpc606_5_976(
      {stage088[21], stage088[22], stage088[23], stage088[24], stage088[25], stage088[26]},
      {stage090[0], stage090[1], stage090[2], stage090[3], stage090[4], stage090[5]},
      {stage092[35], stage091[40], stage090[45], stage089[48], stage088[50]}
   );
   gpc606_5 gpc606_5_977(
      {stage088[27], stage088[28], stage088[29], stage088[30], stage088[31], stage088[32]},
      {stage090[6], stage090[7], stage090[8], stage090[9], stage090[10], stage090[11]},
      {stage092[36], stage091[41], stage090[46], stage089[49], stage088[51]}
   );
   gpc606_5 gpc606_5_978(
      {stage088[33], stage088[34], stage088[35], stage088[36], stage088[37], stage088[38]},
      {stage090[12], stage090[13], stage090[14], stage090[15], stage090[16], stage090[17]},
      {stage092[37], stage091[42], stage090[47], stage089[50], stage088[52]}
   );
   gpc1_1 gpc1_1_979(
      {stage089[25]},
      {stage089[51]}
   );
   gpc1_1 gpc1_1_980(
      {stage089[26]},
      {stage089[52]}
   );
   gpc1_1 gpc1_1_981(
      {stage089[27]},
      {stage089[53]}
   );
   gpc1_1 gpc1_1_982(
      {stage089[28]},
      {stage089[54]}
   );
   gpc1_1 gpc1_1_983(
      {stage089[29]},
      {stage089[55]}
   );
   gpc1_1 gpc1_1_984(
      {stage089[30]},
      {stage089[56]}
   );
   gpc1_1 gpc1_1_985(
      {stage089[31]},
      {stage089[57]}
   );
   gpc623_5 gpc623_5_986(
      {stage089[32], stage089[33], stage089[34]},
      {stage090[18], stage090[19]},
      {stage091[0], stage091[1], stage091[2], stage091[3], stage091[4], stage091[5]},
      {stage093[34], stage092[38], stage091[43], stage090[48], stage089[58]}
   );
   gpc623_5 gpc623_5_987(
      {stage089[35], stage089[36], stage089[37]},
      {stage090[20], stage090[21]},
      {stage091[6], stage091[7], stage091[8], stage091[9], stage091[10], stage091[11]},
      {stage093[35], stage092[39], stage091[44], stage090[49], stage089[59]}
   );
   gpc615_5 gpc615_5_988(
      {stage090[22], stage090[23], stage090[24], stage090[25], stage090[26]},
      {stage091[12]},
      {stage092[0], stage092[1], stage092[2], stage092[3], stage092[4], stage092[5]},
      {stage094[33], stage093[36], stage092[40], stage091[45], stage090[50]}
   );
   gpc615_5 gpc615_5_989(
      {stage090[27], stage090[28], stage090[29], stage090[30], stage090[31]},
      {stage091[13]},
      {stage092[6], stage092[7], stage092[8], stage092[9], stage092[10], stage092[11]},
      {stage094[34], stage093[37], stage092[41], stage091[46], stage090[51]}
   );
   gpc615_5 gpc615_5_990(
      {stage090[32], stage090[33], stage090[34], stage090[35], stage090[36]},
      {stage091[14]},
      {stage092[12], stage092[13], stage092[14], stage092[15], stage092[16], stage092[17]},
      {stage094[35], stage093[38], stage092[42], stage091[47], stage090[52]}
   );
   gpc1_1 gpc1_1_991(
      {stage091[15]},
      {stage091[48]}
   );
   gpc1_1 gpc1_1_992(
      {stage091[16]},
      {stage091[49]}
   );
   gpc1_1 gpc1_1_993(
      {stage091[17]},
      {stage091[50]}
   );
   gpc1_1 gpc1_1_994(
      {stage091[18]},
      {stage091[51]}
   );
   gpc1_1 gpc1_1_995(
      {stage091[19]},
      {stage091[52]}
   );
   gpc1_1 gpc1_1_996(
      {stage091[20]},
      {stage091[53]}
   );
   gpc1_1 gpc1_1_997(
      {stage091[21]},
      {stage091[54]}
   );
   gpc1_1 gpc1_1_998(
      {stage091[22]},
      {stage091[55]}
   );
   gpc1_1 gpc1_1_999(
      {stage091[23]},
      {stage091[56]}
   );
   gpc1_1 gpc1_1_1000(
      {stage091[24]},
      {stage091[57]}
   );
   gpc1_1 gpc1_1_1001(
      {stage091[25]},
      {stage091[58]}
   );
   gpc1_1 gpc1_1_1002(
      {stage091[26]},
      {stage091[59]}
   );
   gpc1_1 gpc1_1_1003(
      {stage091[27]},
      {stage091[60]}
   );
   gpc1_1 gpc1_1_1004(
      {stage091[28]},
      {stage091[61]}
   );
   gpc1_1 gpc1_1_1005(
      {stage091[29]},
      {stage091[62]}
   );
   gpc1_1 gpc1_1_1006(
      {stage091[30]},
      {stage091[63]}
   );
   gpc1_1 gpc1_1_1007(
      {stage091[31]},
      {stage091[64]}
   );
   gpc1_1 gpc1_1_1008(
      {stage091[32]},
      {stage091[65]}
   );
   gpc1_1 gpc1_1_1009(
      {stage091[33]},
      {stage091[66]}
   );
   gpc1_1 gpc1_1_1010(
      {stage091[34]},
      {stage091[67]}
   );
   gpc1_1 gpc1_1_1011(
      {stage091[35]},
      {stage091[68]}
   );
   gpc1_1 gpc1_1_1012(
      {stage092[18]},
      {stage092[43]}
   );
   gpc1_1 gpc1_1_1013(
      {stage092[19]},
      {stage092[44]}
   );
   gpc1_1 gpc1_1_1014(
      {stage092[20]},
      {stage092[45]}
   );
   gpc1_1 gpc1_1_1015(
      {stage092[21]},
      {stage092[46]}
   );
   gpc1_1 gpc1_1_1016(
      {stage092[22]},
      {stage092[47]}
   );
   gpc1_1 gpc1_1_1017(
      {stage092[23]},
      {stage092[48]}
   );
   gpc1_1 gpc1_1_1018(
      {stage092[24]},
      {stage092[49]}
   );
   gpc1_1 gpc1_1_1019(
      {stage092[25]},
      {stage092[50]}
   );
   gpc1_1 gpc1_1_1020(
      {stage092[26]},
      {stage092[51]}
   );
   gpc1_1 gpc1_1_1021(
      {stage092[27]},
      {stage092[52]}
   );
   gpc1_1 gpc1_1_1022(
      {stage092[28]},
      {stage092[53]}
   );
   gpc1_1 gpc1_1_1023(
      {stage092[29]},
      {stage092[54]}
   );
   gpc1_1 gpc1_1_1024(
      {stage092[30]},
      {stage092[55]}
   );
   gpc1_1 gpc1_1_1025(
      {stage092[31]},
      {stage092[56]}
   );
   gpc1_1 gpc1_1_1026(
      {stage092[32]},
      {stage092[57]}
   );
   gpc1_1 gpc1_1_1027(
      {stage092[33]},
      {stage092[58]}
   );
   gpc1_1 gpc1_1_1028(
      {stage092[34]},
      {stage092[59]}
   );
   gpc1_1 gpc1_1_1029(
      {stage093[0]},
      {stage093[39]}
   );
   gpc1_1 gpc1_1_1030(
      {stage093[1]},
      {stage093[40]}
   );
   gpc1_1 gpc1_1_1031(
      {stage093[2]},
      {stage093[41]}
   );
   gpc1_1 gpc1_1_1032(
      {stage093[3]},
      {stage093[42]}
   );
   gpc1_1 gpc1_1_1033(
      {stage093[4]},
      {stage093[43]}
   );
   gpc1_1 gpc1_1_1034(
      {stage093[5]},
      {stage093[44]}
   );
   gpc1_1 gpc1_1_1035(
      {stage093[6]},
      {stage093[45]}
   );
   gpc1_1 gpc1_1_1036(
      {stage093[7]},
      {stage093[46]}
   );
   gpc1_1 gpc1_1_1037(
      {stage093[8]},
      {stage093[47]}
   );
   gpc1_1 gpc1_1_1038(
      {stage093[9]},
      {stage093[48]}
   );
   gpc1_1 gpc1_1_1039(
      {stage093[10]},
      {stage093[49]}
   );
   gpc1_1 gpc1_1_1040(
      {stage093[11]},
      {stage093[50]}
   );
   gpc1_1 gpc1_1_1041(
      {stage093[12]},
      {stage093[51]}
   );
   gpc1_1 gpc1_1_1042(
      {stage093[13]},
      {stage093[52]}
   );
   gpc1_1 gpc1_1_1043(
      {stage093[14]},
      {stage093[53]}
   );
   gpc1_1 gpc1_1_1044(
      {stage093[15]},
      {stage093[54]}
   );
   gpc1_1 gpc1_1_1045(
      {stage093[16]},
      {stage093[55]}
   );
   gpc1_1 gpc1_1_1046(
      {stage093[17]},
      {stage093[56]}
   );
   gpc1_1 gpc1_1_1047(
      {stage093[18]},
      {stage093[57]}
   );
   gpc1_1 gpc1_1_1048(
      {stage093[19]},
      {stage093[58]}
   );
   gpc1_1 gpc1_1_1049(
      {stage093[20]},
      {stage093[59]}
   );
   gpc1_1 gpc1_1_1050(
      {stage093[21]},
      {stage093[60]}
   );
   gpc1_1 gpc1_1_1051(
      {stage093[22]},
      {stage093[61]}
   );
   gpc1_1 gpc1_1_1052(
      {stage093[23]},
      {stage093[62]}
   );
   gpc1_1 gpc1_1_1053(
      {stage093[24]},
      {stage093[63]}
   );
   gpc1_1 gpc1_1_1054(
      {stage093[25]},
      {stage093[64]}
   );
   gpc1_1 gpc1_1_1055(
      {stage093[26]},
      {stage093[65]}
   );
   gpc1_1 gpc1_1_1056(
      {stage093[27]},
      {stage093[66]}
   );
   gpc606_5 gpc606_5_1057(
      {stage093[28], stage093[29], stage093[30], stage093[31], stage093[32], stage093[33]},
      {stage095[0], stage095[1], stage095[2], stage095[3], stage095[4], stage095[5]},
      {stage097[30], stage096[31], stage095[32], stage094[36], stage093[67]}
   );
   gpc1_1 gpc1_1_1058(
      {stage094[0]},
      {stage094[37]}
   );
   gpc1_1 gpc1_1_1059(
      {stage094[1]},
      {stage094[38]}
   );
   gpc1_1 gpc1_1_1060(
      {stage094[2]},
      {stage094[39]}
   );
   gpc1_1 gpc1_1_1061(
      {stage094[3]},
      {stage094[40]}
   );
   gpc1_1 gpc1_1_1062(
      {stage094[4]},
      {stage094[41]}
   );
   gpc1_1 gpc1_1_1063(
      {stage094[5]},
      {stage094[42]}
   );
   gpc1_1 gpc1_1_1064(
      {stage094[6]},
      {stage094[43]}
   );
   gpc1_1 gpc1_1_1065(
      {stage094[7]},
      {stage094[44]}
   );
   gpc1_1 gpc1_1_1066(
      {stage094[8]},
      {stage094[45]}
   );
   gpc1_1 gpc1_1_1067(
      {stage094[9]},
      {stage094[46]}
   );
   gpc1_1 gpc1_1_1068(
      {stage094[10]},
      {stage094[47]}
   );
   gpc1_1 gpc1_1_1069(
      {stage094[11]},
      {stage094[48]}
   );
   gpc1_1 gpc1_1_1070(
      {stage094[12]},
      {stage094[49]}
   );
   gpc1_1 gpc1_1_1071(
      {stage094[13]},
      {stage094[50]}
   );
   gpc1_1 gpc1_1_1072(
      {stage094[14]},
      {stage094[51]}
   );
   gpc606_5 gpc606_5_1073(
      {stage094[15], stage094[16], stage094[17], stage094[18], stage094[19], stage094[20]},
      {stage096[0], stage096[1], stage096[2], stage096[3], stage096[4], stage096[5]},
      {stage098[29], stage097[31], stage096[32], stage095[33], stage094[52]}
   );
   gpc606_5 gpc606_5_1074(
      {stage094[21], stage094[22], stage094[23], stage094[24], stage094[25], stage094[26]},
      {stage096[6], stage096[7], stage096[8], stage096[9], stage096[10], stage096[11]},
      {stage098[30], stage097[32], stage096[33], stage095[34], stage094[53]}
   );
   gpc606_5 gpc606_5_1075(
      {stage094[27], stage094[28], stage094[29], stage094[30], stage094[31], stage094[32]},
      {stage096[12], stage096[13], stage096[14], stage096[15], stage096[16], stage096[17]},
      {stage098[31], stage097[33], stage096[34], stage095[35], stage094[54]}
   );
   gpc1_1 gpc1_1_1076(
      {stage095[6]},
      {stage095[36]}
   );
   gpc1_1 gpc1_1_1077(
      {stage095[7]},
      {stage095[37]}
   );
   gpc1_1 gpc1_1_1078(
      {stage095[8]},
      {stage095[38]}
   );
   gpc1_1 gpc1_1_1079(
      {stage095[9]},
      {stage095[39]}
   );
   gpc1_1 gpc1_1_1080(
      {stage095[10]},
      {stage095[40]}
   );
   gpc1_1 gpc1_1_1081(
      {stage095[11]},
      {stage095[41]}
   );
   gpc1_1 gpc1_1_1082(
      {stage095[12]},
      {stage095[42]}
   );
   gpc1_1 gpc1_1_1083(
      {stage095[13]},
      {stage095[43]}
   );
   gpc1_1 gpc1_1_1084(
      {stage095[14]},
      {stage095[44]}
   );
   gpc1_1 gpc1_1_1085(
      {stage095[15]},
      {stage095[45]}
   );
   gpc1_1 gpc1_1_1086(
      {stage095[16]},
      {stage095[46]}
   );
   gpc1_1 gpc1_1_1087(
      {stage095[17]},
      {stage095[47]}
   );
   gpc1_1 gpc1_1_1088(
      {stage095[18]},
      {stage095[48]}
   );
   gpc1_1 gpc1_1_1089(
      {stage095[19]},
      {stage095[49]}
   );
   gpc1_1 gpc1_1_1090(
      {stage095[20]},
      {stage095[50]}
   );
   gpc1_1 gpc1_1_1091(
      {stage095[21]},
      {stage095[51]}
   );
   gpc1_1 gpc1_1_1092(
      {stage095[22]},
      {stage095[52]}
   );
   gpc1_1 gpc1_1_1093(
      {stage095[23]},
      {stage095[53]}
   );
   gpc1_1 gpc1_1_1094(
      {stage095[24]},
      {stage095[54]}
   );
   gpc1_1 gpc1_1_1095(
      {stage095[25]},
      {stage095[55]}
   );
   gpc606_5 gpc606_5_1096(
      {stage095[26], stage095[27], stage095[28], stage095[29], stage095[30], stage095[31]},
      {stage097[0], stage097[1], stage097[2], stage097[3], stage097[4], stage097[5]},
      {stage099[28], stage098[32], stage097[34], stage096[35], stage095[56]}
   );
   gpc1_1 gpc1_1_1097(
      {stage096[18]},
      {stage096[36]}
   );
   gpc1_1 gpc1_1_1098(
      {stage096[19]},
      {stage096[37]}
   );
   gpc1_1 gpc1_1_1099(
      {stage096[20]},
      {stage096[38]}
   );
   gpc1_1 gpc1_1_1100(
      {stage096[21]},
      {stage096[39]}
   );
   gpc1_1 gpc1_1_1101(
      {stage096[22]},
      {stage096[40]}
   );
   gpc1_1 gpc1_1_1102(
      {stage096[23]},
      {stage096[41]}
   );
   gpc1_1 gpc1_1_1103(
      {stage096[24]},
      {stage096[42]}
   );
   gpc1_1 gpc1_1_1104(
      {stage096[25]},
      {stage096[43]}
   );
   gpc615_5 gpc615_5_1105(
      {stage096[26], stage096[27], stage096[28], stage096[29], stage096[30]},
      {stage097[6]},
      {stage098[0], stage098[1], stage098[2], stage098[3], stage098[4], stage098[5]},
      {stage100[27], stage099[29], stage098[33], stage097[35], stage096[44]}
   );
   gpc1_1 gpc1_1_1106(
      {stage097[7]},
      {stage097[36]}
   );
   gpc1_1 gpc1_1_1107(
      {stage097[8]},
      {stage097[37]}
   );
   gpc1_1 gpc1_1_1108(
      {stage097[9]},
      {stage097[38]}
   );
   gpc615_5 gpc615_5_1109(
      {stage097[10], stage097[11], stage097[12], stage097[13], stage097[14]},
      {stage098[6]},
      {stage099[0], stage099[1], stage099[2], stage099[3], stage099[4], stage099[5]},
      {stage101[26], stage100[28], stage099[30], stage098[34], stage097[39]}
   );
   gpc615_5 gpc615_5_1110(
      {stage097[15], stage097[16], stage097[17], stage097[18], stage097[19]},
      {stage098[7]},
      {stage099[6], stage099[7], stage099[8], stage099[9], stage099[10], stage099[11]},
      {stage101[27], stage100[29], stage099[31], stage098[35], stage097[40]}
   );
   gpc615_5 gpc615_5_1111(
      {stage097[20], stage097[21], stage097[22], stage097[23], stage097[24]},
      {stage098[8]},
      {stage099[12], stage099[13], stage099[14], stage099[15], stage099[16], stage099[17]},
      {stage101[28], stage100[30], stage099[32], stage098[36], stage097[41]}
   );
   gpc615_5 gpc615_5_1112(
      {stage097[25], stage097[26], stage097[27], stage097[28], stage097[29]},
      {stage098[9]},
      {stage099[18], stage099[19], stage099[20], stage099[21], stage099[22], stage099[23]},
      {stage101[29], stage100[31], stage099[33], stage098[37], stage097[42]}
   );
   gpc1_1 gpc1_1_1113(
      {stage098[10]},
      {stage098[38]}
   );
   gpc1_1 gpc1_1_1114(
      {stage098[11]},
      {stage098[39]}
   );
   gpc1_1 gpc1_1_1115(
      {stage098[12]},
      {stage098[40]}
   );
   gpc1_1 gpc1_1_1116(
      {stage098[13]},
      {stage098[41]}
   );
   gpc1_1 gpc1_1_1117(
      {stage098[14]},
      {stage098[42]}
   );
   gpc1_1 gpc1_1_1118(
      {stage098[15]},
      {stage098[43]}
   );
   gpc1_1 gpc1_1_1119(
      {stage098[16]},
      {stage098[44]}
   );
   gpc606_5 gpc606_5_1120(
      {stage098[17], stage098[18], stage098[19], stage098[20], stage098[21], stage098[22]},
      {stage100[0], stage100[1], stage100[2], stage100[3], stage100[4], stage100[5]},
      {stage102[25], stage101[30], stage100[32], stage099[34], stage098[45]}
   );
   gpc606_5 gpc606_5_1121(
      {stage098[23], stage098[24], stage098[25], stage098[26], stage098[27], stage098[28]},
      {stage100[6], stage100[7], stage100[8], stage100[9], stage100[10], stage100[11]},
      {stage102[26], stage101[31], stage100[33], stage099[35], stage098[46]}
   );
   gpc1_1 gpc1_1_1122(
      {stage099[24]},
      {stage099[36]}
   );
   gpc1_1 gpc1_1_1123(
      {stage099[25]},
      {stage099[37]}
   );
   gpc1_1 gpc1_1_1124(
      {stage099[26]},
      {stage099[38]}
   );
   gpc1_1 gpc1_1_1125(
      {stage099[27]},
      {stage099[39]}
   );
   gpc1_1 gpc1_1_1126(
      {stage100[12]},
      {stage100[34]}
   );
   gpc1_1 gpc1_1_1127(
      {stage100[13]},
      {stage100[35]}
   );
   gpc1_1 gpc1_1_1128(
      {stage100[14]},
      {stage100[36]}
   );
   gpc1_1 gpc1_1_1129(
      {stage100[15]},
      {stage100[37]}
   );
   gpc1_1 gpc1_1_1130(
      {stage100[16]},
      {stage100[38]}
   );
   gpc1_1 gpc1_1_1131(
      {stage100[17]},
      {stage100[39]}
   );
   gpc1_1 gpc1_1_1132(
      {stage100[18]},
      {stage100[40]}
   );
   gpc1_1 gpc1_1_1133(
      {stage100[19]},
      {stage100[41]}
   );
   gpc1_1 gpc1_1_1134(
      {stage100[20]},
      {stage100[42]}
   );
   gpc1_1 gpc1_1_1135(
      {stage100[21]},
      {stage100[43]}
   );
   gpc615_5 gpc615_5_1136(
      {stage100[22], stage100[23], stage100[24], stage100[25], stage100[26]},
      {stage101[0]},
      {stage102[0], stage102[1], stage102[2], stage102[3], stage102[4], stage102[5]},
      {stage104[23], stage103[24], stage102[27], stage101[32], stage100[44]}
   );
   gpc1_1 gpc1_1_1137(
      {stage101[1]},
      {stage101[33]}
   );
   gpc1_1 gpc1_1_1138(
      {stage101[2]},
      {stage101[34]}
   );
   gpc7_3 gpc7_3_1139(
      {stage101[3], stage101[4], stage101[5], stage101[6], stage101[7], stage101[8], stage101[9]},
      {stage103[25], stage102[28], stage101[35]}
   );
   gpc606_5 gpc606_5_1140(
      {stage101[10], stage101[11], stage101[12], stage101[13], stage101[14], stage101[15]},
      {stage103[0], stage103[1], stage103[2], stage103[3], stage103[4], stage103[5]},
      {stage105[22], stage104[24], stage103[26], stage102[29], stage101[36]}
   );
   gpc615_5 gpc615_5_1141(
      {stage101[16], stage101[17], stage101[18], stage101[19], stage101[20]},
      {stage102[6]},
      {stage103[6], stage103[7], stage103[8], stage103[9], stage103[10], stage103[11]},
      {stage105[23], stage104[25], stage103[27], stage102[30], stage101[37]}
   );
   gpc615_5 gpc615_5_1142(
      {stage101[21], stage101[22], stage101[23], stage101[24], stage101[25]},
      {stage102[7]},
      {stage103[12], stage103[13], stage103[14], stage103[15], stage103[16], stage103[17]},
      {stage105[24], stage104[26], stage103[28], stage102[31], stage101[38]}
   );
   gpc1_1 gpc1_1_1143(
      {stage102[8]},
      {stage102[32]}
   );
   gpc1_1 gpc1_1_1144(
      {stage102[9]},
      {stage102[33]}
   );
   gpc1_1 gpc1_1_1145(
      {stage102[10]},
      {stage102[34]}
   );
   gpc1_1 gpc1_1_1146(
      {stage102[11]},
      {stage102[35]}
   );
   gpc1_1 gpc1_1_1147(
      {stage102[12]},
      {stage102[36]}
   );
   gpc1_1 gpc1_1_1148(
      {stage102[13]},
      {stage102[37]}
   );
   gpc1_1 gpc1_1_1149(
      {stage102[14]},
      {stage102[38]}
   );
   gpc615_5 gpc615_5_1150(
      {stage102[15], stage102[16], stage102[17], stage102[18], stage102[19]},
      {stage103[18]},
      {stage104[0], stage104[1], stage104[2], stage104[3], stage104[4], stage104[5]},
      {stage106[21], stage105[25], stage104[27], stage103[29], stage102[39]}
   );
   gpc615_5 gpc615_5_1151(
      {stage102[20], stage102[21], stage102[22], stage102[23], stage102[24]},
      {stage103[19]},
      {stage104[6], stage104[7], stage104[8], stage104[9], stage104[10], stage104[11]},
      {stage106[22], stage105[26], stage104[28], stage103[30], stage102[40]}
   );
   gpc1_1 gpc1_1_1152(
      {stage103[20]},
      {stage103[31]}
   );
   gpc1_1 gpc1_1_1153(
      {stage103[21]},
      {stage103[32]}
   );
   gpc1_1 gpc1_1_1154(
      {stage103[22]},
      {stage103[33]}
   );
   gpc1_1 gpc1_1_1155(
      {stage103[23]},
      {stage103[34]}
   );
   gpc1_1 gpc1_1_1156(
      {stage104[12]},
      {stage104[29]}
   );
   gpc615_5 gpc615_5_1157(
      {stage104[13], stage104[14], stage104[15], stage104[16], stage104[17]},
      {stage105[0]},
      {stage106[0], stage106[1], stage106[2], stage106[3], stage106[4], stage106[5]},
      {stage108[19], stage107[20], stage106[23], stage105[27], stage104[30]}
   );
   gpc615_5 gpc615_5_1158(
      {stage104[18], stage104[19], stage104[20], stage104[21], stage104[22]},
      {stage105[1]},
      {stage106[6], stage106[7], stage106[8], stage106[9], stage106[10], stage106[11]},
      {stage108[20], stage107[21], stage106[24], stage105[28], stage104[31]}
   );
   gpc1_1 gpc1_1_1159(
      {stage105[2]},
      {stage105[29]}
   );
   gpc1_1 gpc1_1_1160(
      {stage105[3]},
      {stage105[30]}
   );
   gpc1_1 gpc1_1_1161(
      {stage105[4]},
      {stage105[31]}
   );
   gpc1_1 gpc1_1_1162(
      {stage105[5]},
      {stage105[32]}
   );
   gpc1_1 gpc1_1_1163(
      {stage105[6]},
      {stage105[33]}
   );
   gpc1_1 gpc1_1_1164(
      {stage105[7]},
      {stage105[34]}
   );
   gpc1_1 gpc1_1_1165(
      {stage105[8]},
      {stage105[35]}
   );
   gpc1_1 gpc1_1_1166(
      {stage105[9]},
      {stage105[36]}
   );
   gpc1_1 gpc1_1_1167(
      {stage105[10]},
      {stage105[37]}
   );
   gpc1_1 gpc1_1_1168(
      {stage105[11]},
      {stage105[38]}
   );
   gpc1_1 gpc1_1_1169(
      {stage105[12]},
      {stage105[39]}
   );
   gpc1_1 gpc1_1_1170(
      {stage105[13]},
      {stage105[40]}
   );
   gpc1_1 gpc1_1_1171(
      {stage105[14]},
      {stage105[41]}
   );
   gpc1_1 gpc1_1_1172(
      {stage105[15]},
      {stage105[42]}
   );
   gpc1_1 gpc1_1_1173(
      {stage105[16]},
      {stage105[43]}
   );
   gpc1_1 gpc1_1_1174(
      {stage105[17]},
      {stage105[44]}
   );
   gpc1_1 gpc1_1_1175(
      {stage105[18]},
      {stage105[45]}
   );
   gpc1_1 gpc1_1_1176(
      {stage105[19]},
      {stage105[46]}
   );
   gpc1_1 gpc1_1_1177(
      {stage105[20]},
      {stage105[47]}
   );
   gpc1_1 gpc1_1_1178(
      {stage105[21]},
      {stage105[48]}
   );
   gpc1_1 gpc1_1_1179(
      {stage106[12]},
      {stage106[25]}
   );
   gpc1_1 gpc1_1_1180(
      {stage106[13]},
      {stage106[26]}
   );
   gpc1_1 gpc1_1_1181(
      {stage106[14]},
      {stage106[27]}
   );
   gpc1_1 gpc1_1_1182(
      {stage106[15]},
      {stage106[28]}
   );
   gpc1_1 gpc1_1_1183(
      {stage106[16]},
      {stage106[29]}
   );
   gpc1_1 gpc1_1_1184(
      {stage106[17]},
      {stage106[30]}
   );
   gpc1_1 gpc1_1_1185(
      {stage106[18]},
      {stage106[31]}
   );
   gpc1_1 gpc1_1_1186(
      {stage106[19]},
      {stage106[32]}
   );
   gpc1_1 gpc1_1_1187(
      {stage106[20]},
      {stage106[33]}
   );
   gpc1_1 gpc1_1_1188(
      {stage107[0]},
      {stage107[22]}
   );
   gpc1_1 gpc1_1_1189(
      {stage107[1]},
      {stage107[23]}
   );
   gpc606_5 gpc606_5_1190(
      {stage107[2], stage107[3], stage107[4], stage107[5], stage107[6], stage107[7]},
      {stage109[0], stage109[1], stage109[2], stage109[3], stage109[4], stage109[5]},
      {stage111[16], stage110[17], stage109[18], stage108[21], stage107[24]}
   );
   gpc606_5 gpc606_5_1191(
      {stage107[8], stage107[9], stage107[10], stage107[11], stage107[12], stage107[13]},
      {stage109[6], stage109[7], stage109[8], stage109[9], stage109[10], stage109[11]},
      {stage111[17], stage110[18], stage109[19], stage108[22], stage107[25]}
   );
   gpc606_5 gpc606_5_1192(
      {stage107[14], stage107[15], stage107[16], stage107[17], stage107[18], stage107[19]},
      {stage109[12], stage109[13], stage109[14], stage109[15], stage109[16], stage109[17]},
      {stage111[18], stage110[19], stage109[20], stage108[23], stage107[26]}
   );
   gpc1_1 gpc1_1_1193(
      {stage108[0]},
      {stage108[24]}
   );
   gpc1_1 gpc1_1_1194(
      {stage108[1]},
      {stage108[25]}
   );
   gpc1_1 gpc1_1_1195(
      {stage108[2]},
      {stage108[26]}
   );
   gpc1_1 gpc1_1_1196(
      {stage108[3]},
      {stage108[27]}
   );
   gpc1_1 gpc1_1_1197(
      {stage108[4]},
      {stage108[28]}
   );
   gpc1_1 gpc1_1_1198(
      {stage108[5]},
      {stage108[29]}
   );
   gpc1_1 gpc1_1_1199(
      {stage108[6]},
      {stage108[30]}
   );
   gpc606_5 gpc606_5_1200(
      {stage108[7], stage108[8], stage108[9], stage108[10], stage108[11], stage108[12]},
      {stage110[0], stage110[1], stage110[2], stage110[3], stage110[4], stage110[5]},
      {stage112[15], stage111[19], stage110[20], stage109[21], stage108[31]}
   );
   gpc606_5 gpc606_5_1201(
      {stage108[13], stage108[14], stage108[15], stage108[16], stage108[17], stage108[18]},
      {stage110[6], stage110[7], stage110[8], stage110[9], stage110[10], stage110[11]},
      {stage112[16], stage111[20], stage110[21], stage109[22], stage108[32]}
   );
   gpc1_1 gpc1_1_1202(
      {stage110[12]},
      {stage110[22]}
   );
   gpc1_1 gpc1_1_1203(
      {stage110[13]},
      {stage110[23]}
   );
   gpc1_1 gpc1_1_1204(
      {stage110[14]},
      {stage110[24]}
   );
   gpc1_1 gpc1_1_1205(
      {stage110[15]},
      {stage110[25]}
   );
   gpc1_1 gpc1_1_1206(
      {stage110[16]},
      {stage110[26]}
   );
   gpc1_1 gpc1_1_1207(
      {stage111[0]},
      {stage111[21]}
   );
   gpc1_1 gpc1_1_1208(
      {stage111[1]},
      {stage111[22]}
   );
   gpc1_1 gpc1_1_1209(
      {stage111[2]},
      {stage111[23]}
   );
   gpc1_1 gpc1_1_1210(
      {stage111[3]},
      {stage111[24]}
   );
   gpc1_1 gpc1_1_1211(
      {stage111[4]},
      {stage111[25]}
   );
   gpc1_1 gpc1_1_1212(
      {stage111[5]},
      {stage111[26]}
   );
   gpc1_1 gpc1_1_1213(
      {stage111[6]},
      {stage111[27]}
   );
   gpc1_1 gpc1_1_1214(
      {stage111[7]},
      {stage111[28]}
   );
   gpc1_1 gpc1_1_1215(
      {stage111[8]},
      {stage111[29]}
   );
   gpc1_1 gpc1_1_1216(
      {stage111[9]},
      {stage111[30]}
   );
   gpc606_5 gpc606_5_1217(
      {stage111[10], stage111[11], stage111[12], stage111[13], stage111[14], stage111[15]},
      {stage113[0], stage113[1], stage113[2], stage113[3], stage113[4], stage113[5]},
      {stage115[12], stage114[13], stage113[14], stage112[17], stage111[31]}
   );
   gpc1_1 gpc1_1_1218(
      {stage112[0]},
      {stage112[18]}
   );
   gpc1_1 gpc1_1_1219(
      {stage112[1]},
      {stage112[19]}
   );
   gpc1_1 gpc1_1_1220(
      {stage112[2]},
      {stage112[20]}
   );
   gpc606_5 gpc606_5_1221(
      {stage112[3], stage112[4], stage112[5], stage112[6], stage112[7], stage112[8]},
      {stage114[0], stage114[1], stage114[2], stage114[3], stage114[4], stage114[5]},
      {stage116[11], stage115[13], stage114[14], stage113[15], stage112[21]}
   );
   gpc606_5 gpc606_5_1222(
      {stage112[9], stage112[10], stage112[11], stage112[12], stage112[13], stage112[14]},
      {stage114[6], stage114[7], stage114[8], stage114[9], stage114[10], stage114[11]},
      {stage116[12], stage115[14], stage114[15], stage113[16], stage112[22]}
   );
   gpc1_1 gpc1_1_1223(
      {stage113[6]},
      {stage113[17]}
   );
   gpc1_1 gpc1_1_1224(
      {stage113[7]},
      {stage113[18]}
   );
   gpc1_1 gpc1_1_1225(
      {stage113[8]},
      {stage113[19]}
   );
   gpc1_1 gpc1_1_1226(
      {stage113[9]},
      {stage113[20]}
   );
   gpc1_1 gpc1_1_1227(
      {stage113[10]},
      {stage113[21]}
   );
   gpc1_1 gpc1_1_1228(
      {stage113[11]},
      {stage113[22]}
   );
   gpc1_1 gpc1_1_1229(
      {stage113[12]},
      {stage113[23]}
   );
   gpc1_1 gpc1_1_1230(
      {stage113[13]},
      {stage113[24]}
   );
   gpc1_1 gpc1_1_1231(
      {stage114[12]},
      {stage114[16]}
   );
   gpc1_1 gpc1_1_1232(
      {stage115[0]},
      {stage115[15]}
   );
   gpc1_1 gpc1_1_1233(
      {stage115[1]},
      {stage115[16]}
   );
   gpc1_1 gpc1_1_1234(
      {stage115[2]},
      {stage115[17]}
   );
   gpc1_1 gpc1_1_1235(
      {stage115[3]},
      {stage115[18]}
   );
   gpc1_1 gpc1_1_1236(
      {stage115[4]},
      {stage115[19]}
   );
   gpc1_1 gpc1_1_1237(
      {stage115[5]},
      {stage115[20]}
   );
   gpc1_1 gpc1_1_1238(
      {stage115[6]},
      {stage115[21]}
   );
   gpc1_1 gpc1_1_1239(
      {stage115[7]},
      {stage115[22]}
   );
   gpc1_1 gpc1_1_1240(
      {stage115[8]},
      {stage115[23]}
   );
   gpc1_1 gpc1_1_1241(
      {stage115[9]},
      {stage115[24]}
   );
   gpc1_1 gpc1_1_1242(
      {stage115[10]},
      {stage115[25]}
   );
   gpc1_1 gpc1_1_1243(
      {stage115[11]},
      {stage115[26]}
   );
   gpc1_1 gpc1_1_1244(
      {stage116[0]},
      {stage116[13]}
   );
   gpc1_1 gpc1_1_1245(
      {stage116[1]},
      {stage116[14]}
   );
   gpc1_1 gpc1_1_1246(
      {stage116[2]},
      {stage116[15]}
   );
   gpc1_1 gpc1_1_1247(
      {stage116[3]},
      {stage116[16]}
   );
   gpc1_1 gpc1_1_1248(
      {stage116[4]},
      {stage116[17]}
   );
   gpc1_1 gpc1_1_1249(
      {stage116[5]},
      {stage116[18]}
   );
   gpc1_1 gpc1_1_1250(
      {stage116[6]},
      {stage116[19]}
   );
   gpc1_1 gpc1_1_1251(
      {stage116[7]},
      {stage116[20]}
   );
   gpc1_1 gpc1_1_1252(
      {stage116[8]},
      {stage116[21]}
   );
   gpc1_1 gpc1_1_1253(
      {stage116[9]},
      {stage116[22]}
   );
   gpc1_1 gpc1_1_1254(
      {stage116[10]},
      {stage116[23]}
   );
   gpc1_1 gpc1_1_1255(
      {stage117[0]},
      {stage117[10]}
   );
   gpc1_1 gpc1_1_1256(
      {stage117[1]},
      {stage117[11]}
   );
   gpc1_1 gpc1_1_1257(
      {stage117[2]},
      {stage117[12]}
   );
   gpc1_1 gpc1_1_1258(
      {stage117[3]},
      {stage117[13]}
   );
   gpc1_1 gpc1_1_1259(
      {stage117[4]},
      {stage117[14]}
   );
   gpc1_1 gpc1_1_1260(
      {stage117[5]},
      {stage117[15]}
   );
   gpc1_1 gpc1_1_1261(
      {stage117[6]},
      {stage117[16]}
   );
   gpc1_1 gpc1_1_1262(
      {stage117[7]},
      {stage117[17]}
   );
   gpc1_1 gpc1_1_1263(
      {stage117[8]},
      {stage117[18]}
   );
   gpc1_1 gpc1_1_1264(
      {stage117[9]},
      {stage117[19]}
   );
   gpc1_1 gpc1_1_1265(
      {stage118[0]},
      {stage118[9]}
   );
   gpc1_1 gpc1_1_1266(
      {stage118[1]},
      {stage118[10]}
   );
   gpc1_1 gpc1_1_1267(
      {stage118[2]},
      {stage118[11]}
   );
   gpc606_5 gpc606_5_1268(
      {stage118[3], stage118[4], stage118[5], stage118[6], stage118[7], stage118[8]},
      {stage120[0], stage120[1], stage120[2], stage120[3], stage120[4], stage120[5]},
      {stage122[5], stage121[6], stage120[7], stage119[8], stage118[12]}
   );
   gpc1_1 gpc1_1_1269(
      {stage119[0]},
      {stage119[9]}
   );
   gpc1_1 gpc1_1_1270(
      {stage119[1]},
      {stage119[10]}
   );
   gpc1_1 gpc1_1_1271(
      {stage119[2]},
      {stage119[11]}
   );
   gpc1_1 gpc1_1_1272(
      {stage119[3]},
      {stage119[12]}
   );
   gpc1_1 gpc1_1_1273(
      {stage119[4]},
      {stage119[13]}
   );
   gpc1_1 gpc1_1_1274(
      {stage119[5]},
      {stage119[14]}
   );
   gpc1_1 gpc1_1_1275(
      {stage119[6]},
      {stage119[15]}
   );
   gpc1_1 gpc1_1_1276(
      {stage119[7]},
      {stage119[16]}
   );
   gpc1_1 gpc1_1_1277(
      {stage120[6]},
      {stage120[8]}
   );
   gpc1_1 gpc1_1_1278(
      {stage121[0]},
      {stage121[7]}
   );
   gpc1_1 gpc1_1_1279(
      {stage121[1]},
      {stage121[8]}
   );
   gpc1_1 gpc1_1_1280(
      {stage121[2]},
      {stage121[9]}
   );
   gpc1343_5 gpc1343_5_1281(
      {stage121[3], stage121[4], stage121[5]},
      {stage122[0], stage122[1], stage122[2], stage122[3]},
      {stage123[0], stage123[1], stage123[2]},
      {stage124[0]},
      {stage125[2], stage124[3], stage123[4], stage122[6], stage121[10]}
   );
   gpc1_1 gpc1_1_1282(
      {stage122[4]},
      {stage122[7]}
   );
   gpc1_1 gpc1_1_1283(
      {stage123[3]},
      {stage123[5]}
   );
   gpc1_1 gpc1_1_1284(
      {stage124[1]},
      {stage124[4]}
   );
   gpc1_1 gpc1_1_1285(
      {stage124[2]},
      {stage124[5]}
   );
   gpc1_1 gpc1_1_1286(
      {stage125[0]},
      {stage125[3]}
   );
   gpc1_1 gpc1_1_1287(
      {stage125[1]},
      {stage125[4]}
   );
   gpc1_1 gpc1_1_1288(
      {stage126[0]},
      {stage126[1]}
   );
   gpc1_1 gpc1_1_1289(
      {stage000[1]},
      {stage000[2]}
   );
   gpc1_1 gpc1_1_1290(
      {stage001[2]},
      {stage001[3]}
   );
   gpc1_1 gpc1_1_1291(
      {stage002[3]},
      {stage002[4]}
   );
   gpc1_1 gpc1_1_1292(
      {stage003[4]},
      {stage003[6]}
   );
   gpc1_1 gpc1_1_1293(
      {stage003[5]},
      {stage003[7]}
   );
   gpc615_5 gpc615_5_1294(
      {stage004[5], stage004[6], stage004[7], stage004[8], stage004[9]},
      {stage005[6]},
      {stage006[7], stage006[8], stage006[9], stage006[10], stage006[11], stage006[12]},
      {stage008[14], stage007[16], stage006[14], stage005[13], stage004[10]}
   );
   gpc1_1 gpc1_1_1295(
      {stage005[7]},
      {stage005[14]}
   );
   gpc1_1 gpc1_1_1296(
      {stage005[8]},
      {stage005[15]}
   );
   gpc1_1 gpc1_1_1297(
      {stage005[9]},
      {stage005[16]}
   );
   gpc1_1 gpc1_1_1298(
      {stage005[10]},
      {stage005[17]}
   );
   gpc1_1 gpc1_1_1299(
      {stage005[11]},
      {stage005[18]}
   );
   gpc1_1 gpc1_1_1300(
      {stage005[12]},
      {stage005[19]}
   );
   gpc1_1 gpc1_1_1301(
      {stage006[13]},
      {stage006[15]}
   );
   gpc1_1 gpc1_1_1302(
      {stage007[8]},
      {stage007[17]}
   );
   gpc1_1 gpc1_1_1303(
      {stage007[9]},
      {stage007[18]}
   );
   gpc1_1 gpc1_1_1304(
      {stage007[10]},
      {stage007[19]}
   );
   gpc1_1 gpc1_1_1305(
      {stage007[11]},
      {stage007[20]}
   );
   gpc1_1 gpc1_1_1306(
      {stage007[12]},
      {stage007[21]}
   );
   gpc1_1 gpc1_1_1307(
      {stage007[13]},
      {stage007[22]}
   );
   gpc1_1 gpc1_1_1308(
      {stage007[14]},
      {stage007[23]}
   );
   gpc1_1 gpc1_1_1309(
      {stage007[15]},
      {stage007[24]}
   );
   gpc1_1 gpc1_1_1310(
      {stage008[9]},
      {stage008[15]}
   );
   gpc1_1 gpc1_1_1311(
      {stage008[10]},
      {stage008[16]}
   );
   gpc1_1 gpc1_1_1312(
      {stage008[11]},
      {stage008[17]}
   );
   gpc1_1 gpc1_1_1313(
      {stage008[12]},
      {stage008[18]}
   );
   gpc1_1 gpc1_1_1314(
      {stage008[13]},
      {stage008[19]}
   );
   gpc1_1 gpc1_1_1315(
      {stage009[10]},
      {stage009[20]}
   );
   gpc1_1 gpc1_1_1316(
      {stage009[11]},
      {stage009[21]}
   );
   gpc1_1 gpc1_1_1317(
      {stage009[12]},
      {stage009[22]}
   );
   gpc1_1 gpc1_1_1318(
      {stage009[13]},
      {stage009[23]}
   );
   gpc1_1 gpc1_1_1319(
      {stage009[14]},
      {stage009[24]}
   );
   gpc1_1 gpc1_1_1320(
      {stage009[15]},
      {stage009[25]}
   );
   gpc1_1 gpc1_1_1321(
      {stage009[16]},
      {stage009[26]}
   );
   gpc1_1 gpc1_1_1322(
      {stage009[17]},
      {stage009[27]}
   );
   gpc1_1 gpc1_1_1323(
      {stage009[18]},
      {stage009[28]}
   );
   gpc1_1 gpc1_1_1324(
      {stage009[19]},
      {stage009[29]}
   );
   gpc1_1 gpc1_1_1325(
      {stage010[11]},
      {stage010[13]}
   );
   gpc1_1 gpc1_1_1326(
      {stage010[12]},
      {stage010[14]}
   );
   gpc1_1 gpc1_1_1327(
      {stage011[12]},
      {stage011[25]}
   );
   gpc606_5 gpc606_5_1328(
      {stage011[13], stage011[14], stage011[15], stage011[16], stage011[17], stage011[18]},
      {stage013[14], stage013[15], stage013[16], stage013[17], stage013[18], stage013[19]},
      {stage015[26], stage014[21], stage013[26], stage012[17], stage011[26]}
   );
   gpc606_5 gpc606_5_1329(
      {stage011[19], stage011[20], stage011[21], stage011[22], stage011[23], stage011[24]},
      {stage013[20], stage013[21], stage013[22], stage013[23], stage013[24], stage013[25]},
      {stage015[27], stage014[22], stage013[27], stage012[18], stage011[27]}
   );
   gpc1_1 gpc1_1_1330(
      {stage012[13]},
      {stage012[19]}
   );
   gpc1_1 gpc1_1_1331(
      {stage012[14]},
      {stage012[20]}
   );
   gpc1_1 gpc1_1_1332(
      {stage012[15]},
      {stage012[21]}
   );
   gpc1_1 gpc1_1_1333(
      {stage012[16]},
      {stage012[22]}
   );
   gpc606_5 gpc606_5_1334(
      {1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0},
      {stage015[16], stage015[17], stage015[18], stage015[19], stage015[20], stage015[21]},
      {stage017[34], stage016[26], stage015[28], stage014[23], stage013[28]}
   );
   gpc1_1 gpc1_1_1335(
      {stage014[15]},
      {stage014[24]}
   );
   gpc1_1 gpc1_1_1336(
      {stage014[16]},
      {stage014[25]}
   );
   gpc1_1 gpc1_1_1337(
      {stage014[17]},
      {stage014[26]}
   );
   gpc1_1 gpc1_1_1338(
      {stage014[18]},
      {stage014[27]}
   );
   gpc1_1 gpc1_1_1339(
      {stage014[19]},
      {stage014[28]}
   );
   gpc1_1 gpc1_1_1340(
      {stage014[20]},
      {stage014[29]}
   );
   gpc1_1 gpc1_1_1341(
      {stage015[22]},
      {stage015[29]}
   );
   gpc1_1 gpc1_1_1342(
      {stage015[23]},
      {stage015[30]}
   );
   gpc1_1 gpc1_1_1343(
      {stage015[24]},
      {stage015[31]}
   );
   gpc1_1 gpc1_1_1344(
      {stage015[25]},
      {stage015[32]}
   );
   gpc1_1 gpc1_1_1345(
      {stage016[17]},
      {stage016[27]}
   );
   gpc1_1 gpc1_1_1346(
      {stage016[18]},
      {stage016[28]}
   );
   gpc1_1 gpc1_1_1347(
      {stage016[19]},
      {stage016[29]}
   );
   gpc1406_5 gpc1406_5_1348(
      {stage016[20], stage016[21], stage016[22], stage016[23], stage016[24], stage016[25]},
      {stage018[19], stage018[20], stage018[21], stage018[22]},
      {stage019[20]},
      {stage020[35], stage019[34], stage018[25], stage017[35], stage016[30]}
   );
   gpc1_1 gpc1_1_1349(
      {stage017[18]},
      {stage017[36]}
   );
   gpc1_1 gpc1_1_1350(
      {stage017[19]},
      {stage017[37]}
   );
   gpc1_1 gpc1_1_1351(
      {stage017[20]},
      {stage017[38]}
   );
   gpc1_1 gpc1_1_1352(
      {stage017[21]},
      {stage017[39]}
   );
   gpc1_1 gpc1_1_1353(
      {stage017[22]},
      {stage017[40]}
   );
   gpc1_1 gpc1_1_1354(
      {stage017[23]},
      {stage017[41]}
   );
   gpc1_1 gpc1_1_1355(
      {stage017[24]},
      {stage017[42]}
   );
   gpc1_1 gpc1_1_1356(
      {stage017[25]},
      {stage017[43]}
   );
   gpc1_1 gpc1_1_1357(
      {stage017[26]},
      {stage017[44]}
   );
   gpc1_1 gpc1_1_1358(
      {stage017[27]},
      {stage017[45]}
   );
   gpc1_1 gpc1_1_1359(
      {stage017[28]},
      {stage017[46]}
   );
   gpc1_1 gpc1_1_1360(
      {stage017[29]},
      {stage017[47]}
   );
   gpc1_1 gpc1_1_1361(
      {stage017[30]},
      {stage017[48]}
   );
   gpc1_1 gpc1_1_1362(
      {stage017[31]},
      {stage017[49]}
   );
   gpc1_1 gpc1_1_1363(
      {stage017[32]},
      {stage017[50]}
   );
   gpc1_1 gpc1_1_1364(
      {stage017[33]},
      {stage017[51]}
   );
   gpc1_1 gpc1_1_1365(
      {stage018[23]},
      {stage018[26]}
   );
   gpc1_1 gpc1_1_1366(
      {stage018[24]},
      {stage018[27]}
   );
   gpc1_1 gpc1_1_1367(
      {stage019[21]},
      {stage019[35]}
   );
   gpc1_1 gpc1_1_1368(
      {stage019[22]},
      {stage019[36]}
   );
   gpc1_1 gpc1_1_1369(
      {stage019[23]},
      {stage019[37]}
   );
   gpc1_1 gpc1_1_1370(
      {stage019[24]},
      {stage019[38]}
   );
   gpc1_1 gpc1_1_1371(
      {stage019[25]},
      {stage019[39]}
   );
   gpc1_1 gpc1_1_1372(
      {stage019[26]},
      {stage019[40]}
   );
   gpc1_1 gpc1_1_1373(
      {stage019[27]},
      {stage019[41]}
   );
   gpc1_1 gpc1_1_1374(
      {stage019[28]},
      {stage019[42]}
   );
   gpc1_1 gpc1_1_1375(
      {stage019[29]},
      {stage019[43]}
   );
   gpc1_1 gpc1_1_1376(
      {stage019[30]},
      {stage019[44]}
   );
   gpc1_1 gpc1_1_1377(
      {stage019[31]},
      {stage019[45]}
   );
   gpc1_1 gpc1_1_1378(
      {stage019[32]},
      {stage019[46]}
   );
   gpc1_1 gpc1_1_1379(
      {stage019[33]},
      {stage019[47]}
   );
   gpc1_1 gpc1_1_1380(
      {stage020[21]},
      {stage020[36]}
   );
   gpc1_1 gpc1_1_1381(
      {stage020[22]},
      {stage020[37]}
   );
   gpc1_1 gpc1_1_1382(
      {stage020[23]},
      {stage020[38]}
   );
   gpc1_1 gpc1_1_1383(
      {stage020[24]},
      {stage020[39]}
   );
   gpc1_1 gpc1_1_1384(
      {stage020[25]},
      {stage020[40]}
   );
   gpc1_1 gpc1_1_1385(
      {stage020[26]},
      {stage020[41]}
   );
   gpc1_1 gpc1_1_1386(
      {stage020[27]},
      {stage020[42]}
   );
   gpc1_1 gpc1_1_1387(
      {stage020[28]},
      {stage020[43]}
   );
   gpc1_1 gpc1_1_1388(
      {stage020[29]},
      {stage020[44]}
   );
   gpc615_5 gpc615_5_1389(
      {stage020[30], stage020[31], stage020[32], stage020[33], stage020[34]},
      {stage021[22]},
      {stage022[23], stage022[24], stage022[25], stage022[26], stage022[27], stage022[28]},
      {stage024[32], stage023[45], stage022[42], stage021[32], stage020[45]}
   );
   gpc1_1 gpc1_1_1390(
      {stage021[23]},
      {stage021[33]}
   );
   gpc1_1 gpc1_1_1391(
      {stage021[24]},
      {stage021[34]}
   );
   gpc1_1 gpc1_1_1392(
      {stage021[25]},
      {stage021[35]}
   );
   gpc1_1 gpc1_1_1393(
      {stage021[26]},
      {stage021[36]}
   );
   gpc1_1 gpc1_1_1394(
      {stage021[27]},
      {stage021[37]}
   );
   gpc1_1 gpc1_1_1395(
      {stage021[28]},
      {stage021[38]}
   );
   gpc1_1 gpc1_1_1396(
      {stage021[29]},
      {stage021[39]}
   );
   gpc1_1 gpc1_1_1397(
      {stage021[30]},
      {stage021[40]}
   );
   gpc1_1 gpc1_1_1398(
      {stage021[31]},
      {stage021[41]}
   );
   gpc1_1 gpc1_1_1399(
      {stage022[29]},
      {stage022[43]}
   );
   gpc1_1 gpc1_1_1400(
      {stage022[30]},
      {stage022[44]}
   );
   gpc1_1 gpc1_1_1401(
      {stage022[31]},
      {stage022[45]}
   );
   gpc1_1 gpc1_1_1402(
      {stage022[32]},
      {stage022[46]}
   );
   gpc1_1 gpc1_1_1403(
      {stage022[33]},
      {stage022[47]}
   );
   gpc1_1 gpc1_1_1404(
      {stage022[34]},
      {stage022[48]}
   );
   gpc1_1 gpc1_1_1405(
      {stage022[35]},
      {stage022[49]}
   );
   gpc1_1 gpc1_1_1406(
      {stage022[36]},
      {stage022[50]}
   );
   gpc1_1 gpc1_1_1407(
      {stage022[37]},
      {stage022[51]}
   );
   gpc1_1 gpc1_1_1408(
      {stage022[38]},
      {stage022[52]}
   );
   gpc1_1 gpc1_1_1409(
      {stage022[39]},
      {stage022[53]}
   );
   gpc1_1 gpc1_1_1410(
      {stage022[40]},
      {stage022[54]}
   );
   gpc1_1 gpc1_1_1411(
      {stage022[41]},
      {stage022[55]}
   );
   gpc1_1 gpc1_1_1412(
      {stage023[24]},
      {stage023[46]}
   );
   gpc1_1 gpc1_1_1413(
      {stage023[25]},
      {stage023[47]}
   );
   gpc1_1 gpc1_1_1414(
      {stage023[26]},
      {stage023[48]}
   );
   gpc1_1 gpc1_1_1415(
      {stage023[27]},
      {stage023[49]}
   );
   gpc1_1 gpc1_1_1416(
      {stage023[28]},
      {stage023[50]}
   );
   gpc1_1 gpc1_1_1417(
      {stage023[29]},
      {stage023[51]}
   );
   gpc1_1 gpc1_1_1418(
      {stage023[30]},
      {stage023[52]}
   );
   gpc1_1 gpc1_1_1419(
      {stage023[31]},
      {stage023[53]}
   );
   gpc1_1 gpc1_1_1420(
      {stage023[32]},
      {stage023[54]}
   );
   gpc606_5 gpc606_5_1421(
      {stage023[33], stage023[34], stage023[35], stage023[36], stage023[37], stage023[38]},
      {stage025[26], stage025[27], stage025[28], stage025[29], stage025[30], stage025[31]},
      {stage027[52], stage026[43], stage025[48], stage024[33], stage023[55]}
   );
   gpc606_5 gpc606_5_1422(
      {stage023[39], stage023[40], stage023[41], stage023[42], stage023[43], stage023[44]},
      {stage025[32], stage025[33], stage025[34], stage025[35], stage025[36], stage025[37]},
      {stage027[53], stage026[44], stage025[49], stage024[34], stage023[56]}
   );
   gpc1_1 gpc1_1_1423(
      {stage024[25]},
      {stage024[35]}
   );
   gpc606_5 gpc606_5_1424(
      {stage024[26], stage024[27], stage024[28], stage024[29], stage024[30], stage024[31]},
      {stage026[27], stage026[28], stage026[29], stage026[30], stage026[31], stage026[32]},
      {stage028[41], stage027[54], stage026[45], stage025[50], stage024[36]}
   );
   gpc1_1 gpc1_1_1425(
      {stage025[38]},
      {stage025[51]}
   );
   gpc1_1 gpc1_1_1426(
      {stage025[39]},
      {stage025[52]}
   );
   gpc1_1 gpc1_1_1427(
      {stage025[40]},
      {stage025[53]}
   );
   gpc1_1 gpc1_1_1428(
      {stage025[41]},
      {stage025[54]}
   );
   gpc1_1 gpc1_1_1429(
      {stage025[42]},
      {stage025[55]}
   );
   gpc1_1 gpc1_1_1430(
      {stage025[43]},
      {stage025[56]}
   );
   gpc1_1 gpc1_1_1431(
      {stage025[44]},
      {stage025[57]}
   );
   gpc1_1 gpc1_1_1432(
      {stage025[45]},
      {stage025[58]}
   );
   gpc1_1 gpc1_1_1433(
      {stage025[46]},
      {stage025[59]}
   );
   gpc1_1 gpc1_1_1434(
      {stage025[47]},
      {stage025[60]}
   );
   gpc1_1 gpc1_1_1435(
      {stage026[33]},
      {stage026[46]}
   );
   gpc1_1 gpc1_1_1436(
      {stage026[34]},
      {stage026[47]}
   );
   gpc1_1 gpc1_1_1437(
      {stage026[35]},
      {stage026[48]}
   );
   gpc1_1 gpc1_1_1438(
      {stage026[36]},
      {stage026[49]}
   );
   gpc1_1 gpc1_1_1439(
      {stage026[37]},
      {stage026[50]}
   );
   gpc1_1 gpc1_1_1440(
      {stage026[38]},
      {stage026[51]}
   );
   gpc1_1 gpc1_1_1441(
      {stage026[39]},
      {stage026[52]}
   );
   gpc1_1 gpc1_1_1442(
      {stage026[40]},
      {stage026[53]}
   );
   gpc1_1 gpc1_1_1443(
      {stage026[41]},
      {stage026[54]}
   );
   gpc1_1 gpc1_1_1444(
      {stage026[42]},
      {stage026[55]}
   );
   gpc1_1 gpc1_1_1445(
      {stage027[28]},
      {stage027[55]}
   );
   gpc1_1 gpc1_1_1446(
      {stage027[29]},
      {stage027[56]}
   );
   gpc1_1 gpc1_1_1447(
      {stage027[30]},
      {stage027[57]}
   );
   gpc1_1 gpc1_1_1448(
      {stage027[31]},
      {stage027[58]}
   );
   gpc1_1 gpc1_1_1449(
      {stage027[32]},
      {stage027[59]}
   );
   gpc1_1 gpc1_1_1450(
      {stage027[33]},
      {stage027[60]}
   );
   gpc1_1 gpc1_1_1451(
      {stage027[34]},
      {stage027[61]}
   );
   gpc1_1 gpc1_1_1452(
      {stage027[35]},
      {stage027[62]}
   );
   gpc1_1 gpc1_1_1453(
      {stage027[36]},
      {stage027[63]}
   );
   gpc1_1 gpc1_1_1454(
      {stage027[37]},
      {stage027[64]}
   );
   gpc1_1 gpc1_1_1455(
      {stage027[38]},
      {stage027[65]}
   );
   gpc1_1 gpc1_1_1456(
      {stage027[39]},
      {stage027[66]}
   );
   gpc1_1 gpc1_1_1457(
      {stage027[40]},
      {stage027[67]}
   );
   gpc1_1 gpc1_1_1458(
      {stage027[41]},
      {stage027[68]}
   );
   gpc1_1 gpc1_1_1459(
      {stage027[42]},
      {stage027[69]}
   );
   gpc1_1 gpc1_1_1460(
      {stage027[43]},
      {stage027[70]}
   );
   gpc1_1 gpc1_1_1461(
      {stage027[44]},
      {stage027[71]}
   );
   gpc1_1 gpc1_1_1462(
      {stage027[45]},
      {stage027[72]}
   );
   gpc1_1 gpc1_1_1463(
      {stage027[46]},
      {stage027[73]}
   );
   gpc1_1 gpc1_1_1464(
      {stage027[47]},
      {stage027[74]}
   );
   gpc1_1 gpc1_1_1465(
      {stage027[48]},
      {stage027[75]}
   );
   gpc1_1 gpc1_1_1466(
      {stage027[49]},
      {stage027[76]}
   );
   gpc1_1 gpc1_1_1467(
      {stage027[50]},
      {stage027[77]}
   );
   gpc1_1 gpc1_1_1468(
      {stage027[51]},
      {stage027[78]}
   );
   gpc1_1 gpc1_1_1469(
      {stage028[29]},
      {stage028[42]}
   );
   gpc1_1 gpc1_1_1470(
      {stage028[30]},
      {stage028[43]}
   );
   gpc1_1 gpc1_1_1471(
      {stage028[31]},
      {stage028[44]}
   );
   gpc1_1 gpc1_1_1472(
      {stage028[32]},
      {stage028[45]}
   );
   gpc1_1 gpc1_1_1473(
      {stage028[33]},
      {stage028[46]}
   );
   gpc1_1 gpc1_1_1474(
      {stage028[34]},
      {stage028[47]}
   );
   gpc606_5 gpc606_5_1475(
      {stage028[35], stage028[36], stage028[37], stage028[38], stage028[39], stage028[40]},
      {stage030[31], stage030[32], stage030[33], stage030[34], stage030[35], stage030[36]},
      {stage032[66], stage031[50], stage030[46], stage029[49], stage028[48]}
   );
   gpc1_1 gpc1_1_1476(
      {stage029[30]},
      {stage029[50]}
   );
   gpc1_1 gpc1_1_1477(
      {stage029[31]},
      {stage029[51]}
   );
   gpc1_1 gpc1_1_1478(
      {stage029[32]},
      {stage029[52]}
   );
   gpc1_1 gpc1_1_1479(
      {stage029[33]},
      {stage029[53]}
   );
   gpc1_1 gpc1_1_1480(
      {stage029[34]},
      {stage029[54]}
   );
   gpc1_1 gpc1_1_1481(
      {stage029[35]},
      {stage029[55]}
   );
   gpc1_1 gpc1_1_1482(
      {stage029[36]},
      {stage029[56]}
   );
   gpc1_1 gpc1_1_1483(
      {stage029[37]},
      {stage029[57]}
   );
   gpc1_1 gpc1_1_1484(
      {stage029[38]},
      {stage029[58]}
   );
   gpc615_5 gpc615_5_1485(
      {stage029[39], stage029[40], stage029[41], stage029[42], stage029[43]},
      {stage030[37]},
      {stage031[32], stage031[33], stage031[34], stage031[35], stage031[36], stage031[37]},
      {stage033[43], stage032[67], stage031[51], stage030[47], stage029[59]}
   );
   gpc615_5 gpc615_5_1486(
      {stage029[44], stage029[45], stage029[46], stage029[47], stage029[48]},
      {stage030[38]},
      {stage031[38], stage031[39], stage031[40], stage031[41], stage031[42], stage031[43]},
      {stage033[44], stage032[68], stage031[52], stage030[48], stage029[60]}
   );
   gpc1_1 gpc1_1_1487(
      {stage030[39]},
      {stage030[49]}
   );
   gpc1_1 gpc1_1_1488(
      {stage030[40]},
      {stage030[50]}
   );
   gpc1_1 gpc1_1_1489(
      {stage030[41]},
      {stage030[51]}
   );
   gpc1_1 gpc1_1_1490(
      {stage030[42]},
      {stage030[52]}
   );
   gpc1_1 gpc1_1_1491(
      {stage030[43]},
      {stage030[53]}
   );
   gpc1_1 gpc1_1_1492(
      {stage030[44]},
      {stage030[54]}
   );
   gpc1_1 gpc1_1_1493(
      {stage030[45]},
      {stage030[55]}
   );
   gpc1_1 gpc1_1_1494(
      {stage031[44]},
      {stage031[53]}
   );
   gpc1_1 gpc1_1_1495(
      {stage031[45]},
      {stage031[54]}
   );
   gpc1_1 gpc1_1_1496(
      {stage031[46]},
      {stage031[55]}
   );
   gpc1_1 gpc1_1_1497(
      {stage031[47]},
      {stage031[56]}
   );
   gpc1_1 gpc1_1_1498(
      {stage031[48]},
      {stage031[57]}
   );
   gpc1_1 gpc1_1_1499(
      {stage031[49]},
      {stage031[58]}
   );
   gpc1_1 gpc1_1_1500(
      {stage032[33]},
      {stage032[69]}
   );
   gpc1_1 gpc1_1_1501(
      {stage032[34]},
      {stage032[70]}
   );
   gpc1_1 gpc1_1_1502(
      {stage032[35]},
      {stage032[71]}
   );
   gpc1_1 gpc1_1_1503(
      {stage032[36]},
      {stage032[72]}
   );
   gpc1_1 gpc1_1_1504(
      {stage032[37]},
      {stage032[73]}
   );
   gpc1_1 gpc1_1_1505(
      {stage032[38]},
      {stage032[74]}
   );
   gpc1_1 gpc1_1_1506(
      {stage032[39]},
      {stage032[75]}
   );
   gpc1_1 gpc1_1_1507(
      {stage032[40]},
      {stage032[76]}
   );
   gpc1_1 gpc1_1_1508(
      {stage032[41]},
      {stage032[77]}
   );
   gpc1_1 gpc1_1_1509(
      {stage032[42]},
      {stage032[78]}
   );
   gpc1_1 gpc1_1_1510(
      {stage032[43]},
      {stage032[79]}
   );
   gpc1_1 gpc1_1_1511(
      {stage032[44]},
      {stage032[80]}
   );
   gpc1_1 gpc1_1_1512(
      {stage032[45]},
      {stage032[81]}
   );
   gpc1_1 gpc1_1_1513(
      {stage032[46]},
      {stage032[82]}
   );
   gpc1_1 gpc1_1_1514(
      {stage032[47]},
      {stage032[83]}
   );
   gpc606_5 gpc606_5_1515(
      {stage032[48], stage032[49], stage032[50], stage032[51], stage032[52], stage032[53]},
      {stage034[35], stage034[36], stage034[37], stage034[38], stage034[39], stage034[40]},
      {stage036[49], stage035[50], stage034[58], stage033[45], stage032[84]}
   );
   gpc606_5 gpc606_5_1516(
      {stage032[54], stage032[55], stage032[56], stage032[57], stage032[58], stage032[59]},
      {stage034[41], stage034[42], stage034[43], stage034[44], stage034[45], stage034[46]},
      {stage036[50], stage035[51], stage034[59], stage033[46], stage032[85]}
   );
   gpc606_5 gpc606_5_1517(
      {stage032[60], stage032[61], stage032[62], stage032[63], stage032[64], stage032[65]},
      {stage034[47], stage034[48], stage034[49], stage034[50], stage034[51], stage034[52]},
      {stage036[51], stage035[52], stage034[60], stage033[47], stage032[86]}
   );
   gpc615_5 gpc615_5_1518(
      {stage033[34], stage033[35], stage033[36], stage033[37], stage033[38]},
      {stage034[53]},
      {stage035[36], stage035[37], stage035[38], stage035[39], stage035[40], stage035[41]},
      {stage037[55], stage036[52], stage035[53], stage034[61], stage033[48]}
   );
   gpc615_5 gpc615_5_1519(
      {stage033[39], stage033[40], stage033[41], stage033[42], 1'h0},
      {stage034[54]},
      {stage035[42], stage035[43], stage035[44], stage035[45], stage035[46], stage035[47]},
      {stage037[56], stage036[53], stage035[54], stage034[62], stage033[49]}
   );
   gpc1_1 gpc1_1_1520(
      {stage034[55]},
      {stage034[63]}
   );
   gpc1_1 gpc1_1_1521(
      {stage034[56]},
      {stage034[64]}
   );
   gpc1_1 gpc1_1_1522(
      {stage034[57]},
      {stage034[65]}
   );
   gpc1_1 gpc1_1_1523(
      {stage035[48]},
      {stage035[55]}
   );
   gpc1_1 gpc1_1_1524(
      {stage035[49]},
      {stage035[56]}
   );
   gpc1_1 gpc1_1_1525(
      {stage036[37]},
      {stage036[54]}
   );
   gpc1_1 gpc1_1_1526(
      {stage036[38]},
      {stage036[55]}
   );
   gpc1_1 gpc1_1_1527(
      {stage036[39]},
      {stage036[56]}
   );
   gpc1_1 gpc1_1_1528(
      {stage036[40]},
      {stage036[57]}
   );
   gpc1_1 gpc1_1_1529(
      {stage036[41]},
      {stage036[58]}
   );
   gpc1_1 gpc1_1_1530(
      {stage036[42]},
      {stage036[59]}
   );
   gpc606_5 gpc606_5_1531(
      {stage036[43], stage036[44], stage036[45], stage036[46], stage036[47], stage036[48]},
      {stage038[39], stage038[40], stage038[41], stage038[42], stage038[43], stage038[44]},
      {stage040[56], stage039[56], stage038[64], stage037[57], stage036[60]}
   );
   gpc1_1 gpc1_1_1532(
      {stage037[38]},
      {stage037[58]}
   );
   gpc1_1 gpc1_1_1533(
      {stage037[39]},
      {stage037[59]}
   );
   gpc1_1 gpc1_1_1534(
      {stage037[40]},
      {stage037[60]}
   );
   gpc1_1 gpc1_1_1535(
      {stage037[41]},
      {stage037[61]}
   );
   gpc1_1 gpc1_1_1536(
      {stage037[42]},
      {stage037[62]}
   );
   gpc1_1 gpc1_1_1537(
      {stage037[43]},
      {stage037[63]}
   );
   gpc1_1 gpc1_1_1538(
      {stage037[44]},
      {stage037[64]}
   );
   gpc615_5 gpc615_5_1539(
      {stage037[45], stage037[46], stage037[47], stage037[48], stage037[49]},
      {stage038[45]},
      {stage039[40], stage039[41], stage039[42], stage039[43], stage039[44], stage039[45]},
      {stage041[63], stage040[57], stage039[57], stage038[65], stage037[65]}
   );
   gpc615_5 gpc615_5_1540(
      {stage037[50], stage037[51], stage037[52], stage037[53], stage037[54]},
      {stage038[46]},
      {stage039[46], stage039[47], stage039[48], stage039[49], stage039[50], stage039[51]},
      {stage041[64], stage040[58], stage039[58], stage038[66], stage037[66]}
   );
   gpc1_1 gpc1_1_1541(
      {stage038[47]},
      {stage038[67]}
   );
   gpc1_1 gpc1_1_1542(
      {stage038[48]},
      {stage038[68]}
   );
   gpc1_1 gpc1_1_1543(
      {stage038[49]},
      {stage038[69]}
   );
   gpc1_1 gpc1_1_1544(
      {stage038[50]},
      {stage038[70]}
   );
   gpc1_1 gpc1_1_1545(
      {stage038[51]},
      {stage038[71]}
   );
   gpc1_1 gpc1_1_1546(
      {stage038[52]},
      {stage038[72]}
   );
   gpc1_1 gpc1_1_1547(
      {stage038[53]},
      {stage038[73]}
   );
   gpc1_1 gpc1_1_1548(
      {stage038[54]},
      {stage038[74]}
   );
   gpc1_1 gpc1_1_1549(
      {stage038[55]},
      {stage038[75]}
   );
   gpc1_1 gpc1_1_1550(
      {stage038[56]},
      {stage038[76]}
   );
   gpc1_1 gpc1_1_1551(
      {stage038[57]},
      {stage038[77]}
   );
   gpc1_1 gpc1_1_1552(
      {stage038[58]},
      {stage038[78]}
   );
   gpc1_1 gpc1_1_1553(
      {stage038[59]},
      {stage038[79]}
   );
   gpc1_1 gpc1_1_1554(
      {stage038[60]},
      {stage038[80]}
   );
   gpc1_1 gpc1_1_1555(
      {stage038[61]},
      {stage038[81]}
   );
   gpc1_1 gpc1_1_1556(
      {stage038[62]},
      {stage038[82]}
   );
   gpc1_1 gpc1_1_1557(
      {stage038[63]},
      {stage038[83]}
   );
   gpc615_5 gpc615_5_1558(
      {stage039[52], stage039[53], stage039[54], stage039[55], 1'h0},
      {stage040[41]},
      {stage041[42], stage041[43], stage041[44], stage041[45], stage041[46], stage041[47]},
      {stage043[64], stage042[67], stage041[65], stage040[59], stage039[59]}
   );
   gpc1_1 gpc1_1_1559(
      {stage040[42]},
      {stage040[60]}
   );
   gpc1_1 gpc1_1_1560(
      {stage040[43]},
      {stage040[61]}
   );
   gpc1_1 gpc1_1_1561(
      {stage040[44]},
      {stage040[62]}
   );
   gpc1_1 gpc1_1_1562(
      {stage040[45]},
      {stage040[63]}
   );
   gpc1_1 gpc1_1_1563(
      {stage040[46]},
      {stage040[64]}
   );
   gpc1_1 gpc1_1_1564(
      {stage040[47]},
      {stage040[65]}
   );
   gpc1_1 gpc1_1_1565(
      {stage040[48]},
      {stage040[66]}
   );
   gpc1_1 gpc1_1_1566(
      {stage040[49]},
      {stage040[67]}
   );
   gpc1_1 gpc1_1_1567(
      {stage040[50]},
      {stage040[68]}
   );
   gpc1_1 gpc1_1_1568(
      {stage040[51]},
      {stage040[69]}
   );
   gpc1_1 gpc1_1_1569(
      {stage040[52]},
      {stage040[70]}
   );
   gpc1_1 gpc1_1_1570(
      {stage040[53]},
      {stage040[71]}
   );
   gpc1_1 gpc1_1_1571(
      {stage040[54]},
      {stage040[72]}
   );
   gpc1_1 gpc1_1_1572(
      {stage040[55]},
      {stage040[73]}
   );
   gpc1_1 gpc1_1_1573(
      {stage041[48]},
      {stage041[66]}
   );
   gpc1_1 gpc1_1_1574(
      {stage041[49]},
      {stage041[67]}
   );
   gpc1_1 gpc1_1_1575(
      {stage041[50]},
      {stage041[68]}
   );
   gpc1_1 gpc1_1_1576(
      {stage041[51]},
      {stage041[69]}
   );
   gpc1_1 gpc1_1_1577(
      {stage041[52]},
      {stage041[70]}
   );
   gpc1_1 gpc1_1_1578(
      {stage041[53]},
      {stage041[71]}
   );
   gpc1_1 gpc1_1_1579(
      {stage041[54]},
      {stage041[72]}
   );
   gpc1_1 gpc1_1_1580(
      {stage041[55]},
      {stage041[73]}
   );
   gpc1_1 gpc1_1_1581(
      {stage041[56]},
      {stage041[74]}
   );
   gpc1_1 gpc1_1_1582(
      {stage041[57]},
      {stage041[75]}
   );
   gpc1415_5 gpc1415_5_1583(
      {stage041[58], stage041[59], stage041[60], stage041[61], stage041[62]},
      {stage042[43]},
      {stage043[44], stage043[45], stage043[46], stage043[47]},
      {stage044[45]},
      {stage045[69], stage044[72], stage043[65], stage042[68], stage041[76]}
   );
   gpc1_1 gpc1_1_1584(
      {stage042[44]},
      {stage042[69]}
   );
   gpc1_1 gpc1_1_1585(
      {stage042[45]},
      {stage042[70]}
   );
   gpc1_1 gpc1_1_1586(
      {stage042[46]},
      {stage042[71]}
   );
   gpc1_1 gpc1_1_1587(
      {stage042[47]},
      {stage042[72]}
   );
   gpc1_1 gpc1_1_1588(
      {stage042[48]},
      {stage042[73]}
   );
   gpc1_1 gpc1_1_1589(
      {stage042[49]},
      {stage042[74]}
   );
   gpc1_1 gpc1_1_1590(
      {stage042[50]},
      {stage042[75]}
   );
   gpc606_5 gpc606_5_1591(
      {stage042[51], stage042[52], stage042[53], stage042[54], stage042[55], stage042[56]},
      {stage044[46], stage044[47], stage044[48], stage044[49], stage044[50], stage044[51]},
      {stage046[64], stage045[70], stage044[73], stage043[66], stage042[76]}
   );
   gpc615_5 gpc615_5_1592(
      {stage042[57], stage042[58], stage042[59], stage042[60], stage042[61]},
      {stage043[48]},
      {stage044[52], stage044[53], stage044[54], stage044[55], stage044[56], stage044[57]},
      {stage046[65], stage045[71], stage044[74], stage043[67], stage042[77]}
   );
   gpc615_5 gpc615_5_1593(
      {stage042[62], stage042[63], stage042[64], stage042[65], stage042[66]},
      {stage043[49]},
      {stage044[58], stage044[59], stage044[60], stage044[61], stage044[62], stage044[63]},
      {stage046[66], stage045[72], stage044[75], stage043[68], stage042[78]}
   );
   gpc1_1 gpc1_1_1594(
      {stage043[50]},
      {stage043[69]}
   );
   gpc1_1 gpc1_1_1595(
      {stage043[51]},
      {stage043[70]}
   );
   gpc1_1 gpc1_1_1596(
      {stage043[52]},
      {stage043[71]}
   );
   gpc1_1 gpc1_1_1597(
      {stage043[53]},
      {stage043[72]}
   );
   gpc1_1 gpc1_1_1598(
      {stage043[54]},
      {stage043[73]}
   );
   gpc1_1 gpc1_1_1599(
      {stage043[55]},
      {stage043[74]}
   );
   gpc1_1 gpc1_1_1600(
      {stage043[56]},
      {stage043[75]}
   );
   gpc1_1 gpc1_1_1601(
      {stage043[57]},
      {stage043[76]}
   );
   gpc1_1 gpc1_1_1602(
      {stage043[58]},
      {stage043[77]}
   );
   gpc1_1 gpc1_1_1603(
      {stage043[59]},
      {stage043[78]}
   );
   gpc1_1 gpc1_1_1604(
      {stage043[60]},
      {stage043[79]}
   );
   gpc1_1 gpc1_1_1605(
      {stage043[61]},
      {stage043[80]}
   );
   gpc1_1 gpc1_1_1606(
      {stage043[62]},
      {stage043[81]}
   );
   gpc1_1 gpc1_1_1607(
      {stage043[63]},
      {stage043[82]}
   );
   gpc1_1 gpc1_1_1608(
      {stage044[64]},
      {stage044[76]}
   );
   gpc1_1 gpc1_1_1609(
      {stage044[65]},
      {stage044[77]}
   );
   gpc606_5 gpc606_5_1610(
      {stage044[66], stage044[67], stage044[68], stage044[69], stage044[70], stage044[71]},
      {stage046[47], stage046[48], stage046[49], stage046[50], stage046[51], stage046[52]},
      {stage048[87], stage047[92], stage046[67], stage045[73], stage044[78]}
   );
   gpc606_5 gpc606_5_1611(
      {stage045[46], stage045[47], stage045[48], stage045[49], stage045[50], stage045[51]},
      {stage047[48], stage047[49], stage047[50], stage047[51], stage047[52], stage047[53]},
      {stage049[72], stage048[88], stage047[93], stage046[68], stage045[74]}
   );
   gpc606_5 gpc606_5_1612(
      {stage045[52], stage045[53], stage045[54], stage045[55], stage045[56], stage045[57]},
      {stage047[54], stage047[55], stage047[56], stage047[57], stage047[58], stage047[59]},
      {stage049[73], stage048[89], stage047[94], stage046[69], stage045[75]}
   );
   gpc606_5 gpc606_5_1613(
      {stage045[58], stage045[59], stage045[60], stage045[61], stage045[62], stage045[63]},
      {stage047[60], stage047[61], stage047[62], stage047[63], stage047[64], stage047[65]},
      {stage049[74], stage048[90], stage047[95], stage046[70], stage045[76]}
   );
   gpc615_5 gpc615_5_1614(
      {stage045[64], stage045[65], stage045[66], stage045[67], stage045[68]},
      {stage046[53]},
      {stage047[66], stage047[67], stage047[68], stage047[69], stage047[70], stage047[71]},
      {stage049[75], stage048[91], stage047[96], stage046[71], stage045[77]}
   );
   gpc1_1 gpc1_1_1615(
      {stage046[54]},
      {stage046[72]}
   );
   gpc1_1 gpc1_1_1616(
      {stage046[55]},
      {stage046[73]}
   );
   gpc1_1 gpc1_1_1617(
      {stage046[56]},
      {stage046[74]}
   );
   gpc1_1 gpc1_1_1618(
      {stage046[57]},
      {stage046[75]}
   );
   gpc1_1 gpc1_1_1619(
      {stage046[58]},
      {stage046[76]}
   );
   gpc1_1 gpc1_1_1620(
      {stage046[59]},
      {stage046[77]}
   );
   gpc1_1 gpc1_1_1621(
      {stage046[60]},
      {stage046[78]}
   );
   gpc1_1 gpc1_1_1622(
      {stage046[61]},
      {stage046[79]}
   );
   gpc1_1 gpc1_1_1623(
      {stage046[62]},
      {stage046[80]}
   );
   gpc1_1 gpc1_1_1624(
      {stage046[63]},
      {stage046[81]}
   );
   gpc1_1 gpc1_1_1625(
      {stage047[72]},
      {stage047[97]}
   );
   gpc1_1 gpc1_1_1626(
      {stage047[73]},
      {stage047[98]}
   );
   gpc606_5 gpc606_5_1627(
      {stage047[74], stage047[75], stage047[76], stage047[77], stage047[78], stage047[79]},
      {stage049[50], stage049[51], stage049[52], stage049[53], stage049[54], stage049[55]},
      {stage051[68], stage050[76], stage049[76], stage048[92], stage047[99]}
   );
   gpc606_5 gpc606_5_1628(
      {stage047[80], stage047[81], stage047[82], stage047[83], stage047[84], stage047[85]},
      {stage049[56], stage049[57], stage049[58], stage049[59], stage049[60], stage049[61]},
      {stage051[69], stage050[77], stage049[77], stage048[93], stage047[100]}
   );
   gpc606_5 gpc606_5_1629(
      {stage047[86], stage047[87], stage047[88], stage047[89], stage047[90], stage047[91]},
      {stage049[62], stage049[63], stage049[64], stage049[65], stage049[66], stage049[67]},
      {stage051[70], stage050[78], stage049[78], stage048[94], stage047[101]}
   );
   gpc1_1 gpc1_1_1630(
      {stage048[49]},
      {stage048[95]}
   );
   gpc1_1 gpc1_1_1631(
      {stage048[50]},
      {stage048[96]}
   );
   gpc1_1 gpc1_1_1632(
      {stage048[51]},
      {stage048[97]}
   );
   gpc1_1 gpc1_1_1633(
      {stage048[52]},
      {stage048[98]}
   );
   gpc1_1 gpc1_1_1634(
      {stage048[53]},
      {stage048[99]}
   );
   gpc1_1 gpc1_1_1635(
      {stage048[54]},
      {stage048[100]}
   );
   gpc1_1 gpc1_1_1636(
      {stage048[55]},
      {stage048[101]}
   );
   gpc1_1 gpc1_1_1637(
      {stage048[56]},
      {stage048[102]}
   );
   gpc1_1 gpc1_1_1638(
      {stage048[57]},
      {stage048[103]}
   );
   gpc1_1 gpc1_1_1639(
      {stage048[58]},
      {stage048[104]}
   );
   gpc1_1 gpc1_1_1640(
      {stage048[59]},
      {stage048[105]}
   );
   gpc1_1 gpc1_1_1641(
      {stage048[60]},
      {stage048[106]}
   );
   gpc1_1 gpc1_1_1642(
      {stage048[61]},
      {stage048[107]}
   );
   gpc1_1 gpc1_1_1643(
      {stage048[62]},
      {stage048[108]}
   );
   gpc1_1 gpc1_1_1644(
      {stage048[63]},
      {stage048[109]}
   );
   gpc1_1 gpc1_1_1645(
      {stage048[64]},
      {stage048[110]}
   );
   gpc1_1 gpc1_1_1646(
      {stage048[65]},
      {stage048[111]}
   );
   gpc1_1 gpc1_1_1647(
      {stage048[66]},
      {stage048[112]}
   );
   gpc1_1 gpc1_1_1648(
      {stage048[67]},
      {stage048[113]}
   );
   gpc1_1 gpc1_1_1649(
      {stage048[68]},
      {stage048[114]}
   );
   gpc606_5 gpc606_5_1650(
      {stage048[69], stage048[70], stage048[71], stage048[72], stage048[73], stage048[74]},
      {stage050[51], stage050[52], stage050[53], stage050[54], stage050[55], stage050[56]},
      {stage052[84], stage051[71], stage050[79], stage049[79], stage048[115]}
   );
   gpc606_5 gpc606_5_1651(
      {stage048[75], stage048[76], stage048[77], stage048[78], stage048[79], stage048[80]},
      {stage050[57], stage050[58], stage050[59], stage050[60], stage050[61], stage050[62]},
      {stage052[85], stage051[72], stage050[80], stage049[80], stage048[116]}
   );
   gpc606_5 gpc606_5_1652(
      {stage048[81], stage048[82], stage048[83], stage048[84], stage048[85], stage048[86]},
      {stage050[63], stage050[64], stage050[65], stage050[66], stage050[67], stage050[68]},
      {stage052[86], stage051[73], stage050[81], stage049[81], stage048[117]}
   );
   gpc1_1 gpc1_1_1653(
      {stage049[68]},
      {stage049[82]}
   );
   gpc1_1 gpc1_1_1654(
      {stage049[69]},
      {stage049[83]}
   );
   gpc1_1 gpc1_1_1655(
      {stage049[70]},
      {stage049[84]}
   );
   gpc1_1 gpc1_1_1656(
      {stage049[71]},
      {stage049[85]}
   );
   gpc1_1 gpc1_1_1657(
      {stage050[69]},
      {stage050[82]}
   );
   gpc1_1 gpc1_1_1658(
      {stage050[70]},
      {stage050[83]}
   );
   gpc1_1 gpc1_1_1659(
      {stage050[71]},
      {stage050[84]}
   );
   gpc1_1 gpc1_1_1660(
      {stage050[72]},
      {stage050[85]}
   );
   gpc1_1 gpc1_1_1661(
      {stage050[73]},
      {stage050[86]}
   );
   gpc1_1 gpc1_1_1662(
      {stage050[74]},
      {stage050[87]}
   );
   gpc1_1 gpc1_1_1663(
      {stage050[75]},
      {stage050[88]}
   );
   gpc1_1 gpc1_1_1664(
      {stage051[52]},
      {stage051[74]}
   );
   gpc615_5 gpc615_5_1665(
      {stage051[53], stage051[54], stage051[55], stage051[56], stage051[57]},
      {stage052[53]},
      {stage053[54], stage053[55], stage053[56], stage053[57], stage053[58], stage053[59]},
      {stage055[84], stage054[100], stage053[101], stage052[87], stage051[75]}
   );
   gpc615_5 gpc615_5_1666(
      {stage051[58], stage051[59], stage051[60], stage051[61], stage051[62]},
      {stage052[54]},
      {stage053[60], stage053[61], stage053[62], stage053[63], stage053[64], stage053[65]},
      {stage055[85], stage054[101], stage053[102], stage052[88], stage051[76]}
   );
   gpc615_5 gpc615_5_1667(
      {stage051[63], stage051[64], stage051[65], stage051[66], stage051[67]},
      {stage052[55]},
      {stage053[66], stage053[67], stage053[68], stage053[69], stage053[70], stage053[71]},
      {stage055[86], stage054[102], stage053[103], stage052[89], stage051[77]}
   );
   gpc1_1 gpc1_1_1668(
      {stage052[56]},
      {stage052[90]}
   );
   gpc1_1 gpc1_1_1669(
      {stage052[57]},
      {stage052[91]}
   );
   gpc1_1 gpc1_1_1670(
      {stage052[58]},
      {stage052[92]}
   );
   gpc615_5 gpc615_5_1671(
      {stage052[59], stage052[60], stage052[61], stage052[62], stage052[63]},
      {stage053[72]},
      {stage054[55], stage054[56], stage054[57], stage054[58], stage054[59], stage054[60]},
      {stage056[75], stage055[87], stage054[103], stage053[104], stage052[93]}
   );
   gpc615_5 gpc615_5_1672(
      {stage052[64], stage052[65], stage052[66], stage052[67], stage052[68]},
      {stage053[73]},
      {stage054[61], stage054[62], stage054[63], stage054[64], stage054[65], stage054[66]},
      {stage056[76], stage055[88], stage054[104], stage053[105], stage052[94]}
   );
   gpc615_5 gpc615_5_1673(
      {stage052[69], stage052[70], stage052[71], stage052[72], stage052[73]},
      {stage053[74]},
      {stage054[67], stage054[68], stage054[69], stage054[70], stage054[71], stage054[72]},
      {stage056[77], stage055[89], stage054[105], stage053[106], stage052[95]}
   );
   gpc615_5 gpc615_5_1674(
      {stage052[74], stage052[75], stage052[76], stage052[77], stage052[78]},
      {stage053[75]},
      {stage054[73], stage054[74], stage054[75], stage054[76], stage054[77], stage054[78]},
      {stage056[78], stage055[90], stage054[106], stage053[107], stage052[96]}
   );
   gpc615_5 gpc615_5_1675(
      {stage052[79], stage052[80], stage052[81], stage052[82], stage052[83]},
      {stage053[76]},
      {stage054[79], stage054[80], stage054[81], stage054[82], stage054[83], stage054[84]},
      {stage056[79], stage055[91], stage054[107], stage053[108], stage052[97]}
   );
   gpc1_1 gpc1_1_1676(
      {stage053[77]},
      {stage053[109]}
   );
   gpc1_1 gpc1_1_1677(
      {stage053[78]},
      {stage053[110]}
   );
   gpc1_1 gpc1_1_1678(
      {stage053[79]},
      {stage053[111]}
   );
   gpc1_1 gpc1_1_1679(
      {stage053[80]},
      {stage053[112]}
   );
   gpc1_1 gpc1_1_1680(
      {stage053[81]},
      {stage053[113]}
   );
   gpc1_1 gpc1_1_1681(
      {stage053[82]},
      {stage053[114]}
   );
   gpc1_1 gpc1_1_1682(
      {stage053[83]},
      {stage053[115]}
   );
   gpc1_1 gpc1_1_1683(
      {stage053[84]},
      {stage053[116]}
   );
   gpc1_1 gpc1_1_1684(
      {stage053[85]},
      {stage053[117]}
   );
   gpc1_1 gpc1_1_1685(
      {stage053[86]},
      {stage053[118]}
   );
   gpc1_1 gpc1_1_1686(
      {stage053[87]},
      {stage053[119]}
   );
   gpc1_1 gpc1_1_1687(
      {stage053[88]},
      {stage053[120]}
   );
   gpc615_5 gpc615_5_1688(
      {stage053[89], stage053[90], stage053[91], stage053[92], stage053[93]},
      {stage054[85]},
      {stage055[56], stage055[57], stage055[58], stage055[59], stage055[60], stage055[61]},
      {stage057[79], stage056[80], stage055[92], stage054[108], stage053[121]}
   );
   gpc207_4 gpc207_4_1689(
      {stage053[94], stage053[95], stage053[96], stage053[97], stage053[98], stage053[99], stage053[100]},
      {stage055[62], stage055[63]},
      {stage056[81], stage055[93], stage054[109], stage053[122]}
   );
   gpc1_1 gpc1_1_1690(
      {stage054[86]},
      {stage054[110]}
   );
   gpc1_1 gpc1_1_1691(
      {stage054[87]},
      {stage054[111]}
   );
   gpc1_1 gpc1_1_1692(
      {stage054[88]},
      {stage054[112]}
   );
   gpc1_1 gpc1_1_1693(
      {stage054[89]},
      {stage054[113]}
   );
   gpc615_5 gpc615_5_1694(
      {stage054[90], stage054[91], stage054[92], stage054[93], stage054[94]},
      {stage055[64]},
      {stage056[57], stage056[58], stage056[59], stage056[60], stage056[61], stage056[62]},
      {stage058[83], stage057[80], stage056[82], stage055[94], stage054[114]}
   );
   gpc615_5 gpc615_5_1695(
      {stage054[95], stage054[96], stage054[97], stage054[98], stage054[99]},
      {stage055[65]},
      {stage056[63], stage056[64], stage056[65], stage056[66], stage056[67], stage056[68]},
      {stage058[84], stage057[81], stage056[83], stage055[95], stage054[115]}
   );
   gpc1_1 gpc1_1_1696(
      {stage055[66]},
      {stage055[96]}
   );
   gpc1_1 gpc1_1_1697(
      {stage055[67]},
      {stage055[97]}
   );
   gpc1_1 gpc1_1_1698(
      {stage055[68]},
      {stage055[98]}
   );
   gpc1_1 gpc1_1_1699(
      {stage055[69]},
      {stage055[99]}
   );
   gpc1_1 gpc1_1_1700(
      {stage055[70]},
      {stage055[100]}
   );
   gpc1_1 gpc1_1_1701(
      {stage055[71]},
      {stage055[101]}
   );
   gpc606_5 gpc606_5_1702(
      {stage055[72], stage055[73], stage055[74], stage055[75], stage055[76], stage055[77]},
      {stage057[58], stage057[59], stage057[60], stage057[61], stage057[62], stage057[63]},
      {stage059[91], stage058[85], stage057[82], stage056[84], stage055[102]}
   );
   gpc606_5 gpc606_5_1703(
      {stage055[78], stage055[79], stage055[80], stage055[81], stage055[82], stage055[83]},
      {stage057[64], stage057[65], stage057[66], stage057[67], stage057[68], stage057[69]},
      {stage059[92], stage058[86], stage057[83], stage056[85], stage055[103]}
   );
   gpc606_5 gpc606_5_1704(
      {stage056[69], stage056[70], stage056[71], stage056[72], stage056[73], stage056[74]},
      {stage058[59], stage058[60], stage058[61], stage058[62], stage058[63], stage058[64]},
      {stage060[85], stage059[93], stage058[87], stage057[84], stage056[86]}
   );
   gpc1_1 gpc1_1_1705(
      {stage057[70]},
      {stage057[85]}
   );
   gpc1_1 gpc1_1_1706(
      {stage057[71]},
      {stage057[86]}
   );
   gpc1_1 gpc1_1_1707(
      {stage057[72]},
      {stage057[87]}
   );
   gpc606_5 gpc606_5_1708(
      {stage057[73], stage057[74], stage057[75], stage057[76], stage057[77], stage057[78]},
      {stage059[60], stage059[61], stage059[62], stage059[63], stage059[64], stage059[65]},
      {stage061[103], stage060[86], stage059[94], stage058[88], stage057[88]}
   );
   gpc1_1 gpc1_1_1709(
      {stage058[65]},
      {stage058[89]}
   );
   gpc1_1 gpc1_1_1710(
      {stage058[66]},
      {stage058[90]}
   );
   gpc1_1 gpc1_1_1711(
      {stage058[67]},
      {stage058[91]}
   );
   gpc615_5 gpc615_5_1712(
      {stage058[68], stage058[69], stage058[70], stage058[71], stage058[72]},
      {stage059[66]},
      {stage060[61], stage060[62], stage060[63], stage060[64], stage060[65], stage060[66]},
      {stage062[102], stage061[104], stage060[87], stage059[95], stage058[92]}
   );
   gpc615_5 gpc615_5_1713(
      {stage058[73], stage058[74], stage058[75], stage058[76], stage058[77]},
      {stage059[67]},
      {stage060[67], stage060[68], stage060[69], stage060[70], stage060[71], stage060[72]},
      {stage062[103], stage061[105], stage060[88], stage059[96], stage058[93]}
   );
   gpc2135_5 gpc2135_5_1714(
      {stage058[78], stage058[79], stage058[80], stage058[81], stage058[82]},
      {stage059[68], stage059[69], stage059[70]},
      {stage060[73]},
      {stage061[62], stage061[63]},
      {stage062[104], stage061[106], stage060[89], stage059[97], stage058[94]}
   );
   gpc1_1 gpc1_1_1715(
      {stage059[71]},
      {stage059[98]}
   );
   gpc1_1 gpc1_1_1716(
      {stage059[72]},
      {stage059[99]}
   );
   gpc606_5 gpc606_5_1717(
      {stage059[73], stage059[74], stage059[75], stage059[76], stage059[77], stage059[78]},
      {stage061[64], stage061[65], stage061[66], stage061[67], stage061[68], stage061[69]},
      {stage063[104], stage062[105], stage061[107], stage060[90], stage059[100]}
   );
   gpc606_5 gpc606_5_1718(
      {stage059[79], stage059[80], stage059[81], stage059[82], stage059[83], stage059[84]},
      {stage061[70], stage061[71], stage061[72], stage061[73], stage061[74], stage061[75]},
      {stage063[105], stage062[106], stage061[108], stage060[91], stage059[101]}
   );
   gpc606_5 gpc606_5_1719(
      {stage059[85], stage059[86], stage059[87], stage059[88], stage059[89], stage059[90]},
      {stage061[76], stage061[77], stage061[78], stage061[79], stage061[80], stage061[81]},
      {stage063[106], stage062[107], stage061[109], stage060[92], stage059[102]}
   );
   gpc1_1 gpc1_1_1720(
      {stage060[74]},
      {stage060[93]}
   );
   gpc1_1 gpc1_1_1721(
      {stage060[75]},
      {stage060[94]}
   );
   gpc1_1 gpc1_1_1722(
      {stage060[76]},
      {stage060[95]}
   );
   gpc1_1 gpc1_1_1723(
      {stage060[77]},
      {stage060[96]}
   );
   gpc1_1 gpc1_1_1724(
      {stage060[78]},
      {stage060[97]}
   );
   gpc606_5 gpc606_5_1725(
      {stage060[79], stage060[80], stage060[81], stage060[82], stage060[83], stage060[84]},
      {stage062[63], stage062[64], stage062[65], stage062[66], stage062[67], stage062[68]},
      {stage064[97], stage063[107], stage062[108], stage061[110], stage060[98]}
   );
   gpc1_1 gpc1_1_1726(
      {stage061[82]},
      {stage061[111]}
   );
   gpc1_1 gpc1_1_1727(
      {stage061[83]},
      {stage061[112]}
   );
   gpc1_1 gpc1_1_1728(
      {stage061[84]},
      {stage061[113]}
   );
   gpc1_1 gpc1_1_1729(
      {stage061[85]},
      {stage061[114]}
   );
   gpc1_1 gpc1_1_1730(
      {stage061[86]},
      {stage061[115]}
   );
   gpc1_1 gpc1_1_1731(
      {stage061[87]},
      {stage061[116]}
   );
   gpc615_5 gpc615_5_1732(
      {stage061[88], stage061[89], stage061[90], stage061[91], stage061[92]},
      {stage062[69]},
      {stage063[64], stage063[65], stage063[66], stage063[67], stage063[68], stage063[69]},
      {stage065[91], stage064[98], stage063[108], stage062[109], stage061[117]}
   );
   gpc615_5 gpc615_5_1733(
      {stage061[93], stage061[94], stage061[95], stage061[96], stage061[97]},
      {stage062[70]},
      {stage063[70], stage063[71], stage063[72], stage063[73], stage063[74], stage063[75]},
      {stage065[92], stage064[99], stage063[109], stage062[110], stage061[118]}
   );
   gpc615_5 gpc615_5_1734(
      {stage061[98], stage061[99], stage061[100], stage061[101], stage061[102]},
      {stage062[71]},
      {stage063[76], stage063[77], stage063[78], stage063[79], stage063[80], stage063[81]},
      {stage065[93], stage064[100], stage063[110], stage062[111], stage061[119]}
   );
   gpc1_1 gpc1_1_1735(
      {stage062[72]},
      {stage062[112]}
   );
   gpc1_1 gpc1_1_1736(
      {stage062[73]},
      {stage062[113]}
   );
   gpc1_1 gpc1_1_1737(
      {stage062[74]},
      {stage062[114]}
   );
   gpc1_1 gpc1_1_1738(
      {stage062[75]},
      {stage062[115]}
   );
   gpc1_1 gpc1_1_1739(
      {stage062[76]},
      {stage062[116]}
   );
   gpc1_1 gpc1_1_1740(
      {stage062[77]},
      {stage062[117]}
   );
   gpc1_1 gpc1_1_1741(
      {stage062[78]},
      {stage062[118]}
   );
   gpc1_1 gpc1_1_1742(
      {stage062[79]},
      {stage062[119]}
   );
   gpc1_1 gpc1_1_1743(
      {stage062[80]},
      {stage062[120]}
   );
   gpc1_1 gpc1_1_1744(
      {stage062[81]},
      {stage062[121]}
   );
   gpc615_5 gpc615_5_1745(
      {stage062[82], stage062[83], stage062[84], stage062[85], stage062[86]},
      {stage063[82]},
      {stage064[63], stage064[64], stage064[65], stage064[66], stage064[67], stage064[68]},
      {stage066[85], stage065[94], stage064[101], stage063[111], stage062[122]}
   );
   gpc615_5 gpc615_5_1746(
      {stage062[87], stage062[88], stage062[89], stage062[90], stage062[91]},
      {stage063[83]},
      {stage064[69], stage064[70], stage064[71], stage064[72], stage064[73], stage064[74]},
      {stage066[86], stage065[95], stage064[102], stage063[112], stage062[123]}
   );
   gpc615_5 gpc615_5_1747(
      {stage062[92], stage062[93], stage062[94], stage062[95], stage062[96]},
      {stage063[84]},
      {stage064[75], stage064[76], stage064[77], stage064[78], stage064[79], stage064[80]},
      {stage066[87], stage065[96], stage064[103], stage063[113], stage062[124]}
   );
   gpc615_5 gpc615_5_1748(
      {stage062[97], stage062[98], stage062[99], stage062[100], stage062[101]},
      {stage063[85]},
      {stage064[81], stage064[82], stage064[83], stage064[84], stage064[85], stage064[86]},
      {stage066[88], stage065[97], stage064[104], stage063[114], stage062[125]}
   );
   gpc1_1 gpc1_1_1749(
      {stage063[86]},
      {stage063[115]}
   );
   gpc1_1 gpc1_1_1750(
      {stage063[87]},
      {stage063[116]}
   );
   gpc1_1 gpc1_1_1751(
      {stage063[88]},
      {stage063[117]}
   );
   gpc1_1 gpc1_1_1752(
      {stage063[89]},
      {stage063[118]}
   );
   gpc1_1 gpc1_1_1753(
      {stage063[90]},
      {stage063[119]}
   );
   gpc1_1 gpc1_1_1754(
      {stage063[91]},
      {stage063[120]}
   );
   gpc1_1 gpc1_1_1755(
      {stage063[92]},
      {stage063[121]}
   );
   gpc1_1 gpc1_1_1756(
      {stage063[93]},
      {stage063[122]}
   );
   gpc1_1 gpc1_1_1757(
      {stage063[94]},
      {stage063[123]}
   );
   gpc1_1 gpc1_1_1758(
      {stage063[95]},
      {stage063[124]}
   );
   gpc1_1 gpc1_1_1759(
      {stage063[96]},
      {stage063[125]}
   );
   gpc1_1 gpc1_1_1760(
      {stage063[97]},
      {stage063[126]}
   );
   gpc1_1 gpc1_1_1761(
      {stage063[98]},
      {stage063[127]}
   );
   gpc615_5 gpc615_5_1762(
      {stage063[99], stage063[100], stage063[101], stage063[102], stage063[103]},
      {stage064[87]},
      {stage065[62], stage065[63], stage065[64], stage065[65], stage065[66], stage065[67]},
      {stage067[103], stage066[89], stage065[98], stage064[105], stage063[128]}
   );
   gpc615_5 gpc615_5_1763(
      {stage064[88], stage064[89], stage064[90], stage064[91], stage064[92]},
      {stage065[68]},
      {stage066[61], stage066[62], stage066[63], stage066[64], stage066[65], stage066[66]},
      {stage068[85], stage067[104], stage066[90], stage065[99], stage064[106]}
   );
   gpc615_5 gpc615_5_1764(
      {stage064[93], stage064[94], stage064[95], stage064[96], 1'h0},
      {stage065[69]},
      {stage066[67], stage066[68], stage066[69], stage066[70], stage066[71], stage066[72]},
      {stage068[86], stage067[105], stage066[91], stage065[100], stage064[107]}
   );
   gpc1_1 gpc1_1_1765(
      {stage065[70]},
      {stage065[101]}
   );
   gpc1_1 gpc1_1_1766(
      {stage065[71]},
      {stage065[102]}
   );
   gpc1_1 gpc1_1_1767(
      {stage065[72]},
      {stage065[103]}
   );
   gpc1_1 gpc1_1_1768(
      {stage065[73]},
      {stage065[104]}
   );
   gpc1_1 gpc1_1_1769(
      {stage065[74]},
      {stage065[105]}
   );
   gpc1_1 gpc1_1_1770(
      {stage065[75]},
      {stage065[106]}
   );
   gpc1_1 gpc1_1_1771(
      {stage065[76]},
      {stage065[107]}
   );
   gpc1_1 gpc1_1_1772(
      {stage065[77]},
      {stage065[108]}
   );
   gpc1_1 gpc1_1_1773(
      {stage065[78]},
      {stage065[109]}
   );
   gpc1_1 gpc1_1_1774(
      {stage065[79]},
      {stage065[110]}
   );
   gpc1_1 gpc1_1_1775(
      {stage065[80]},
      {stage065[111]}
   );
   gpc1_1 gpc1_1_1776(
      {stage065[81]},
      {stage065[112]}
   );
   gpc1_1 gpc1_1_1777(
      {stage065[82]},
      {stage065[113]}
   );
   gpc623_5 gpc623_5_1778(
      {stage065[83], stage065[84], stage065[85]},
      {stage066[73], stage066[74]},
      {stage067[60], stage067[61], stage067[62], stage067[63], stage067[64], stage067[65]},
      {stage069[92], stage068[87], stage067[106], stage066[92], stage065[114]}
   );
   gpc615_5 gpc615_5_1779(
      {stage065[86], stage065[87], stage065[88], stage065[89], stage065[90]},
      {stage066[75]},
      {stage067[66], stage067[67], stage067[68], stage067[69], stage067[70], stage067[71]},
      {stage069[93], stage068[88], stage067[107], stage066[93], stage065[115]}
   );
   gpc1_1 gpc1_1_1780(
      {stage066[76]},
      {stage066[94]}
   );
   gpc1_1 gpc1_1_1781(
      {stage066[77]},
      {stage066[95]}
   );
   gpc1_1 gpc1_1_1782(
      {stage066[78]},
      {stage066[96]}
   );
   gpc1_1 gpc1_1_1783(
      {stage066[79]},
      {stage066[97]}
   );
   gpc615_5 gpc615_5_1784(
      {stage066[80], stage066[81], stage066[82], stage066[83], stage066[84]},
      {stage067[72]},
      {stage068[59], stage068[60], stage068[61], stage068[62], stage068[63], stage068[64]},
      {stage070[90], stage069[94], stage068[89], stage067[108], stage066[98]}
   );
   gpc1_1 gpc1_1_1785(
      {stage067[73]},
      {stage067[109]}
   );
   gpc606_5 gpc606_5_1786(
      {stage067[74], stage067[75], stage067[76], stage067[77], stage067[78], stage067[79]},
      {stage069[58], stage069[59], stage069[60], stage069[61], stage069[62], stage069[63]},
      {stage071[80], stage070[91], stage069[95], stage068[90], stage067[110]}
   );
   gpc606_5 gpc606_5_1787(
      {stage067[80], stage067[81], stage067[82], stage067[83], stage067[84], stage067[85]},
      {stage069[64], stage069[65], stage069[66], stage069[67], stage069[68], stage069[69]},
      {stage071[81], stage070[92], stage069[96], stage068[91], stage067[111]}
   );
   gpc606_5 gpc606_5_1788(
      {stage067[86], stage067[87], stage067[88], stage067[89], stage067[90], stage067[91]},
      {stage069[70], stage069[71], stage069[72], stage069[73], stage069[74], stage069[75]},
      {stage071[82], stage070[93], stage069[97], stage068[92], stage067[112]}
   );
   gpc606_5 gpc606_5_1789(
      {stage067[92], stage067[93], stage067[94], stage067[95], stage067[96], stage067[97]},
      {stage069[76], stage069[77], stage069[78], stage069[79], stage069[80], stage069[81]},
      {stage071[83], stage070[94], stage069[98], stage068[93], stage067[113]}
   );
   gpc615_5 gpc615_5_1790(
      {stage067[98], stage067[99], stage067[100], stage067[101], stage067[102]},
      {stage068[65]},
      {stage069[82], stage069[83], stage069[84], stage069[85], stage069[86], stage069[87]},
      {stage071[84], stage070[95], stage069[99], stage068[94], stage067[114]}
   );
   gpc1_1 gpc1_1_1791(
      {stage068[66]},
      {stage068[95]}
   );
   gpc606_5 gpc606_5_1792(
      {stage068[67], stage068[68], stage068[69], stage068[70], stage068[71], stage068[72]},
      {stage070[57], stage070[58], stage070[59], stage070[60], stage070[61], stage070[62]},
      {stage072[83], stage071[85], stage070[96], stage069[100], stage068[96]}
   );
   gpc606_5 gpc606_5_1793(
      {stage068[73], stage068[74], stage068[75], stage068[76], stage068[77], stage068[78]},
      {stage070[63], stage070[64], stage070[65], stage070[66], stage070[67], stage070[68]},
      {stage072[84], stage071[86], stage070[97], stage069[101], stage068[97]}
   );
   gpc606_5 gpc606_5_1794(
      {stage068[79], stage068[80], stage068[81], stage068[82], stage068[83], stage068[84]},
      {stage070[69], stage070[70], stage070[71], stage070[72], stage070[73], stage070[74]},
      {stage072[85], stage071[87], stage070[98], stage069[102], stage068[98]}
   );
   gpc1_1 gpc1_1_1795(
      {stage069[88]},
      {stage069[103]}
   );
   gpc1_1 gpc1_1_1796(
      {stage069[89]},
      {stage069[104]}
   );
   gpc1_1 gpc1_1_1797(
      {stage069[90]},
      {stage069[105]}
   );
   gpc1_1 gpc1_1_1798(
      {stage069[91]},
      {stage069[106]}
   );
   gpc615_5 gpc615_5_1799(
      {stage070[75], stage070[76], stage070[77], stage070[78], stage070[79]},
      {stage071[56]},
      {stage072[55], stage072[56], stage072[57], stage072[58], stage072[59], stage072[60]},
      {stage074[81], stage073[84], stage072[86], stage071[88], stage070[99]}
   );
   gpc615_5 gpc615_5_1800(
      {stage070[80], stage070[81], stage070[82], stage070[83], stage070[84]},
      {stage071[57]},
      {stage072[61], stage072[62], stage072[63], stage072[64], stage072[65], stage072[66]},
      {stage074[82], stage073[85], stage072[87], stage071[89], stage070[100]}
   );
   gpc615_5 gpc615_5_1801(
      {stage070[85], stage070[86], stage070[87], stage070[88], stage070[89]},
      {stage071[58]},
      {stage072[67], stage072[68], stage072[69], stage072[70], stage072[71], stage072[72]},
      {stage074[83], stage073[86], stage072[88], stage071[90], stage070[101]}
   );
   gpc1_1 gpc1_1_1802(
      {stage071[59]},
      {stage071[91]}
   );
   gpc1_1 gpc1_1_1803(
      {stage071[60]},
      {stage071[92]}
   );
   gpc1_1 gpc1_1_1804(
      {stage071[61]},
      {stage071[93]}
   );
   gpc1_1 gpc1_1_1805(
      {stage071[62]},
      {stage071[94]}
   );
   gpc1_1 gpc1_1_1806(
      {stage071[63]},
      {stage071[95]}
   );
   gpc1_1 gpc1_1_1807(
      {stage071[64]},
      {stage071[96]}
   );
   gpc615_5 gpc615_5_1808(
      {stage071[65], stage071[66], stage071[67], stage071[68], stage071[69]},
      {stage072[73]},
      {stage073[54], stage073[55], stage073[56], stage073[57], stage073[58], stage073[59]},
      {stage075[78], stage074[84], stage073[87], stage072[89], stage071[97]}
   );
   gpc615_5 gpc615_5_1809(
      {stage071[70], stage071[71], stage071[72], stage071[73], stage071[74]},
      {stage072[74]},
      {stage073[60], stage073[61], stage073[62], stage073[63], stage073[64], stage073[65]},
      {stage075[79], stage074[85], stage073[88], stage072[90], stage071[98]}
   );
   gpc615_5 gpc615_5_1810(
      {stage071[75], stage071[76], stage071[77], stage071[78], stage071[79]},
      {stage072[75]},
      {stage073[66], stage073[67], stage073[68], stage073[69], stage073[70], stage073[71]},
      {stage075[80], stage074[86], stage073[89], stage072[91], stage071[99]}
   );
   gpc1_1 gpc1_1_1811(
      {stage072[76]},
      {stage072[92]}
   );
   gpc1_1 gpc1_1_1812(
      {stage072[77]},
      {stage072[93]}
   );
   gpc1_1 gpc1_1_1813(
      {stage072[78]},
      {stage072[94]}
   );
   gpc1_1 gpc1_1_1814(
      {stage072[79]},
      {stage072[95]}
   );
   gpc1_1 gpc1_1_1815(
      {stage072[80]},
      {stage072[96]}
   );
   gpc1_1 gpc1_1_1816(
      {stage072[81]},
      {stage072[97]}
   );
   gpc1_1 gpc1_1_1817(
      {stage072[82]},
      {stage072[98]}
   );
   gpc606_5 gpc606_5_1818(
      {stage073[72], stage073[73], stage073[74], stage073[75], stage073[76], stage073[77]},
      {stage075[52], stage075[53], stage075[54], stage075[55], stage075[56], stage075[57]},
      {stage077[75], stage076[73], stage075[81], stage074[87], stage073[90]}
   );
   gpc606_5 gpc606_5_1819(
      {stage073[78], stage073[79], stage073[80], stage073[81], stage073[82], stage073[83]},
      {stage075[58], stage075[59], stage075[60], stage075[61], stage075[62], stage075[63]},
      {stage077[76], stage076[74], stage075[82], stage074[88], stage073[91]}
   );
   gpc1_1 gpc1_1_1820(
      {stage074[53]},
      {stage074[89]}
   );
   gpc1_1 gpc1_1_1821(
      {stage074[54]},
      {stage074[90]}
   );
   gpc1_1 gpc1_1_1822(
      {stage074[55]},
      {stage074[91]}
   );
   gpc1_1 gpc1_1_1823(
      {stage074[56]},
      {stage074[92]}
   );
   gpc1_1 gpc1_1_1824(
      {stage074[57]},
      {stage074[93]}
   );
   gpc1_1 gpc1_1_1825(
      {stage074[58]},
      {stage074[94]}
   );
   gpc1_1 gpc1_1_1826(
      {stage074[59]},
      {stage074[95]}
   );
   gpc1_1 gpc1_1_1827(
      {stage074[60]},
      {stage074[96]}
   );
   gpc1_1 gpc1_1_1828(
      {stage074[61]},
      {stage074[97]}
   );
   gpc1_1 gpc1_1_1829(
      {stage074[62]},
      {stage074[98]}
   );
   gpc1_1 gpc1_1_1830(
      {stage074[63]},
      {stage074[99]}
   );
   gpc1_1 gpc1_1_1831(
      {stage074[64]},
      {stage074[100]}
   );
   gpc1_1 gpc1_1_1832(
      {stage074[65]},
      {stage074[101]}
   );
   gpc615_5 gpc615_5_1833(
      {stage074[66], stage074[67], stage074[68], stage074[69], stage074[70]},
      {stage075[64]},
      {stage076[51], stage076[52], stage076[53], stage076[54], stage076[55], stage076[56]},
      {stage078[71], stage077[77], stage076[75], stage075[83], stage074[102]}
   );
   gpc615_5 gpc615_5_1834(
      {stage074[71], stage074[72], stage074[73], stage074[74], stage074[75]},
      {stage075[65]},
      {stage076[57], stage076[58], stage076[59], stage076[60], stage076[61], stage076[62]},
      {stage078[72], stage077[78], stage076[76], stage075[84], stage074[103]}
   );
   gpc615_5 gpc615_5_1835(
      {stage074[76], stage074[77], stage074[78], stage074[79], stage074[80]},
      {stage075[66]},
      {stage076[63], stage076[64], stage076[65], stage076[66], stage076[67], stage076[68]},
      {stage078[73], stage077[79], stage076[77], stage075[85], stage074[104]}
   );
   gpc606_5 gpc606_5_1836(
      {stage075[67], stage075[68], stage075[69], stage075[70], stage075[71], stage075[72]},
      {stage077[50], stage077[51], stage077[52], stage077[53], stage077[54], stage077[55]},
      {stage079[85], stage078[74], stage077[80], stage076[78], stage075[86]}
   );
   gpc606_5 gpc606_5_1837(
      {stage075[73], stage075[74], stage075[75], stage075[76], stage075[77], 1'h0},
      {stage077[56], stage077[57], stage077[58], stage077[59], stage077[60], stage077[61]},
      {stage079[86], stage078[75], stage077[81], stage076[79], stage075[87]}
   );
   gpc1_1 gpc1_1_1838(
      {stage076[69]},
      {stage076[80]}
   );
   gpc1_1 gpc1_1_1839(
      {stage076[70]},
      {stage076[81]}
   );
   gpc1_1 gpc1_1_1840(
      {stage076[71]},
      {stage076[82]}
   );
   gpc1_1 gpc1_1_1841(
      {stage076[72]},
      {stage076[83]}
   );
   gpc1_1 gpc1_1_1842(
      {stage077[62]},
      {stage077[82]}
   );
   gpc1_1 gpc1_1_1843(
      {stage077[63]},
      {stage077[83]}
   );
   gpc1_1 gpc1_1_1844(
      {stage077[64]},
      {stage077[84]}
   );
   gpc1_1 gpc1_1_1845(
      {stage077[65]},
      {stage077[85]}
   );
   gpc1_1 gpc1_1_1846(
      {stage077[66]},
      {stage077[86]}
   );
   gpc1_1 gpc1_1_1847(
      {stage077[67]},
      {stage077[87]}
   );
   gpc1_1 gpc1_1_1848(
      {stage077[68]},
      {stage077[88]}
   );
   gpc606_5 gpc606_5_1849(
      {stage077[69], stage077[70], stage077[71], stage077[72], stage077[73], stage077[74]},
      {stage079[48], stage079[49], stage079[50], stage079[51], stage079[52], stage079[53]},
      {stage081[75], stage080[71], stage079[87], stage078[76], stage077[89]}
   );
   gpc1_1 gpc1_1_1850(
      {stage078[49]},
      {stage078[77]}
   );
   gpc1_1 gpc1_1_1851(
      {stage078[50]},
      {stage078[78]}
   );
   gpc1_1 gpc1_1_1852(
      {stage078[51]},
      {stage078[79]}
   );
   gpc1_1 gpc1_1_1853(
      {stage078[52]},
      {stage078[80]}
   );
   gpc1_1 gpc1_1_1854(
      {stage078[53]},
      {stage078[81]}
   );
   gpc1_1 gpc1_1_1855(
      {stage078[54]},
      {stage078[82]}
   );
   gpc1_1 gpc1_1_1856(
      {stage078[55]},
      {stage078[83]}
   );
   gpc1_1 gpc1_1_1857(
      {stage078[56]},
      {stage078[84]}
   );
   gpc1_1 gpc1_1_1858(
      {stage078[57]},
      {stage078[85]}
   );
   gpc1_1 gpc1_1_1859(
      {stage078[58]},
      {stage078[86]}
   );
   gpc606_5 gpc606_5_1860(
      {stage078[59], stage078[60], stage078[61], stage078[62], stage078[63], stage078[64]},
      {stage080[47], stage080[48], stage080[49], stage080[50], stage080[51], stage080[52]},
      {stage082[66], stage081[76], stage080[72], stage079[88], stage078[87]}
   );
   gpc606_5 gpc606_5_1861(
      {stage078[65], stage078[66], stage078[67], stage078[68], stage078[69], stage078[70]},
      {stage080[53], stage080[54], stage080[55], stage080[56], stage080[57], stage080[58]},
      {stage082[67], stage081[77], stage080[73], stage079[89], stage078[88]}
   );
   gpc1_1 gpc1_1_1862(
      {stage079[54]},
      {stage079[90]}
   );
   gpc1_1 gpc1_1_1863(
      {stage079[55]},
      {stage079[91]}
   );
   gpc1_1 gpc1_1_1864(
      {stage079[56]},
      {stage079[92]}
   );
   gpc1_1 gpc1_1_1865(
      {stage079[57]},
      {stage079[93]}
   );
   gpc1_1 gpc1_1_1866(
      {stage079[58]},
      {stage079[94]}
   );
   gpc1_1 gpc1_1_1867(
      {stage079[59]},
      {stage079[95]}
   );
   gpc1_1 gpc1_1_1868(
      {stage079[60]},
      {stage079[96]}
   );
   gpc606_5 gpc606_5_1869(
      {stage079[61], stage079[62], stage079[63], stage079[64], stage079[65], stage079[66]},
      {stage081[46], stage081[47], stage081[48], stage081[49], stage081[50], stage081[51]},
      {stage083[63], stage082[68], stage081[78], stage080[74], stage079[97]}
   );
   gpc606_5 gpc606_5_1870(
      {stage079[67], stage079[68], stage079[69], stage079[70], stage079[71], stage079[72]},
      {stage081[52], stage081[53], stage081[54], stage081[55], stage081[56], stage081[57]},
      {stage083[64], stage082[69], stage081[79], stage080[75], stage079[98]}
   );
   gpc606_5 gpc606_5_1871(
      {stage079[73], stage079[74], stage079[75], stage079[76], stage079[77], stage079[78]},
      {stage081[58], stage081[59], stage081[60], stage081[61], stage081[62], stage081[63]},
      {stage083[65], stage082[70], stage081[80], stage080[76], stage079[99]}
   );
   gpc606_5 gpc606_5_1872(
      {stage079[79], stage079[80], stage079[81], stage079[82], stage079[83], stage079[84]},
      {stage081[64], stage081[65], stage081[66], stage081[67], stage081[68], stage081[69]},
      {stage083[66], stage082[71], stage081[81], stage080[77], stage079[100]}
   );
   gpc1_1 gpc1_1_1873(
      {stage080[59]},
      {stage080[78]}
   );
   gpc1_1 gpc1_1_1874(
      {stage080[60]},
      {stage080[79]}
   );
   gpc1_1 gpc1_1_1875(
      {stage080[61]},
      {stage080[80]}
   );
   gpc1_1 gpc1_1_1876(
      {stage080[62]},
      {stage080[81]}
   );
   gpc1_1 gpc1_1_1877(
      {stage080[63]},
      {stage080[82]}
   );
   gpc1_1 gpc1_1_1878(
      {stage080[64]},
      {stage080[83]}
   );
   gpc606_5 gpc606_5_1879(
      {stage080[65], stage080[66], stage080[67], stage080[68], stage080[69], stage080[70]},
      {stage082[45], stage082[46], stage082[47], stage082[48], stage082[49], stage082[50]},
      {stage084[74], stage083[67], stage082[72], stage081[82], stage080[84]}
   );
   gpc1415_5 gpc1415_5_1880(
      {stage081[70], stage081[71], stage081[72], stage081[73], stage081[74]},
      {stage082[51]},
      {stage083[44], stage083[45], stage083[46], stage083[47]},
      {stage084[43]},
      {stage085[68], stage084[75], stage083[68], stage082[73], stage081[83]}
   );
   gpc1_1 gpc1_1_1881(
      {stage082[52]},
      {stage082[74]}
   );
   gpc1_1 gpc1_1_1882(
      {stage082[53]},
      {stage082[75]}
   );
   gpc606_5 gpc606_5_1883(
      {stage082[54], stage082[55], stage082[56], stage082[57], stage082[58], stage082[59]},
      {stage084[44], stage084[45], stage084[46], stage084[47], stage084[48], stage084[49]},
      {stage086[66], stage085[69], stage084[76], stage083[69], stage082[76]}
   );
   gpc606_5 gpc606_5_1884(
      {stage082[60], stage082[61], stage082[62], stage082[63], stage082[64], stage082[65]},
      {stage084[50], stage084[51], stage084[52], stage084[53], stage084[54], stage084[55]},
      {stage086[67], stage085[70], stage084[77], stage083[70], stage082[77]}
   );
   gpc615_5 gpc615_5_1885(
      {stage083[48], stage083[49], stage083[50], stage083[51], stage083[52]},
      {stage084[56]},
      {stage085[42], stage085[43], stage085[44], stage085[45], stage085[46], stage085[47]},
      {stage087[54], stage086[68], stage085[71], stage084[78], stage083[71]}
   );
   gpc615_5 gpc615_5_1886(
      {stage083[53], stage083[54], stage083[55], stage083[56], stage083[57]},
      {stage084[57]},
      {stage085[48], stage085[49], stage085[50], stage085[51], stage085[52], stage085[53]},
      {stage087[55], stage086[69], stage085[72], stage084[79], stage083[72]}
   );
   gpc615_5 gpc615_5_1887(
      {stage083[58], stage083[59], stage083[60], stage083[61], stage083[62]},
      {stage084[58]},
      {stage085[54], stage085[55], stage085[56], stage085[57], stage085[58], stage085[59]},
      {stage087[56], stage086[70], stage085[73], stage084[80], stage083[73]}
   );
   gpc7_3 gpc7_3_1888(
      {stage084[59], stage084[60], stage084[61], stage084[62], stage084[63], stage084[64], stage084[65]},
      {stage086[71], stage085[74], stage084[81]}
   );
   gpc615_5 gpc615_5_1889(
      {stage084[66], stage084[67], stage084[68], stage084[69], stage084[70]},
      {stage085[60]},
      {stage086[41], stage086[42], stage086[43], stage086[44], stage086[45], stage086[46]},
      {stage088[53], stage087[57], stage086[72], stage085[75], stage084[82]}
   );
   gpc615_5 gpc615_5_1890(
      {stage084[71], stage084[72], stage084[73], 1'h0, 1'h0},
      {stage085[61]},
      {stage086[47], stage086[48], stage086[49], stage086[50], stage086[51], stage086[52]},
      {stage088[54], stage087[58], stage086[73], stage085[76], stage084[83]}
   );
   gpc1_1 gpc1_1_1891(
      {stage085[62]},
      {stage085[77]}
   );
   gpc1_1 gpc1_1_1892(
      {stage085[63]},
      {stage085[78]}
   );
   gpc1_1 gpc1_1_1893(
      {stage085[64]},
      {stage085[79]}
   );
   gpc623_5 gpc623_5_1894(
      {stage085[65], stage085[66], stage085[67]},
      {stage086[53], stage086[54]},
      {stage087[40], stage087[41], stage087[42], stage087[43], stage087[44], stage087[45]},
      {stage089[60], stage088[55], stage087[59], stage086[74], stage085[80]}
   );
   gpc1_1 gpc1_1_1895(
      {stage086[55]},
      {stage086[75]}
   );
   gpc1_1 gpc1_1_1896(
      {stage086[56]},
      {stage086[76]}
   );
   gpc1_1 gpc1_1_1897(
      {stage086[57]},
      {stage086[77]}
   );
   gpc1_1 gpc1_1_1898(
      {stage086[58]},
      {stage086[78]}
   );
   gpc1_1 gpc1_1_1899(
      {stage086[59]},
      {stage086[79]}
   );
   gpc606_5 gpc606_5_1900(
      {stage086[60], stage086[61], stage086[62], stage086[63], stage086[64], stage086[65]},
      {stage088[39], stage088[40], stage088[41], stage088[42], stage088[43], stage088[44]},
      {stage090[53], stage089[61], stage088[56], stage087[60], stage086[80]}
   );
   gpc1_1 gpc1_1_1901(
      {stage087[46]},
      {stage087[61]}
   );
   gpc1_1 gpc1_1_1902(
      {stage087[47]},
      {stage087[62]}
   );
   gpc606_5 gpc606_5_1903(
      {stage087[48], stage087[49], stage087[50], stage087[51], stage087[52], stage087[53]},
      {stage089[38], stage089[39], stage089[40], stage089[41], stage089[42], stage089[43]},
      {stage091[69], stage090[54], stage089[62], stage088[57], stage087[63]}
   );
   gpc1_1 gpc1_1_1904(
      {stage088[45]},
      {stage088[58]}
   );
   gpc1_1 gpc1_1_1905(
      {stage088[46]},
      {stage088[59]}
   );
   gpc1_1 gpc1_1_1906(
      {stage088[47]},
      {stage088[60]}
   );
   gpc1_1 gpc1_1_1907(
      {stage088[48]},
      {stage088[61]}
   );
   gpc1_1 gpc1_1_1908(
      {stage088[49]},
      {stage088[62]}
   );
   gpc1_1 gpc1_1_1909(
      {stage088[50]},
      {stage088[63]}
   );
   gpc1_1 gpc1_1_1910(
      {stage088[51]},
      {stage088[64]}
   );
   gpc1_1 gpc1_1_1911(
      {stage088[52]},
      {stage088[65]}
   );
   gpc1_1 gpc1_1_1912(
      {stage089[44]},
      {stage089[63]}
   );
   gpc1_1 gpc1_1_1913(
      {stage089[45]},
      {stage089[64]}
   );
   gpc1_1 gpc1_1_1914(
      {stage089[46]},
      {stage089[65]}
   );
   gpc1_1 gpc1_1_1915(
      {stage089[47]},
      {stage089[66]}
   );
   gpc1_1 gpc1_1_1916(
      {stage089[48]},
      {stage089[67]}
   );
   gpc1_1 gpc1_1_1917(
      {stage089[49]},
      {stage089[68]}
   );
   gpc615_5 gpc615_5_1918(
      {stage089[50], stage089[51], stage089[52], stage089[53], stage089[54]},
      {stage090[37]},
      {stage091[36], stage091[37], stage091[38], stage091[39], stage091[40], stage091[41]},
      {stage093[68], stage092[60], stage091[70], stage090[55], stage089[69]}
   );
   gpc615_5 gpc615_5_1919(
      {stage089[55], stage089[56], stage089[57], stage089[58], stage089[59]},
      {stage090[38]},
      {stage091[42], stage091[43], stage091[44], stage091[45], stage091[46], stage091[47]},
      {stage093[69], stage092[61], stage091[71], stage090[56], stage089[70]}
   );
   gpc1_1 gpc1_1_1920(
      {stage090[39]},
      {stage090[57]}
   );
   gpc1_1 gpc1_1_1921(
      {stage090[40]},
      {stage090[58]}
   );
   gpc1_1 gpc1_1_1922(
      {stage090[41]},
      {stage090[59]}
   );
   gpc1_1 gpc1_1_1923(
      {stage090[42]},
      {stage090[60]}
   );
   gpc1_1 gpc1_1_1924(
      {stage090[43]},
      {stage090[61]}
   );
   gpc1_1 gpc1_1_1925(
      {stage090[44]},
      {stage090[62]}
   );
   gpc1_1 gpc1_1_1926(
      {stage090[45]},
      {stage090[63]}
   );
   gpc1_1 gpc1_1_1927(
      {stage090[46]},
      {stage090[64]}
   );
   gpc1_1 gpc1_1_1928(
      {stage090[47]},
      {stage090[65]}
   );
   gpc615_5 gpc615_5_1929(
      {stage090[48], stage090[49], stage090[50], stage090[51], stage090[52]},
      {stage091[48]},
      {stage092[35], stage092[36], stage092[37], stage092[38], stage092[39], stage092[40]},
      {stage094[55], stage093[70], stage092[62], stage091[72], stage090[66]}
   );
   gpc1_1 gpc1_1_1930(
      {stage091[49]},
      {stage091[73]}
   );
   gpc1_1 gpc1_1_1931(
      {stage091[50]},
      {stage091[74]}
   );
   gpc1_1 gpc1_1_1932(
      {stage091[51]},
      {stage091[75]}
   );
   gpc1_1 gpc1_1_1933(
      {stage091[52]},
      {stage091[76]}
   );
   gpc606_5 gpc606_5_1934(
      {stage091[53], stage091[54], stage091[55], stage091[56], stage091[57], stage091[58]},
      {stage093[34], stage093[35], stage093[36], stage093[37], stage093[38], stage093[39]},
      {stage095[57], stage094[56], stage093[71], stage092[63], stage091[77]}
   );
   gpc615_5 gpc615_5_1935(
      {stage091[59], stage091[60], stage091[61], stage091[62], stage091[63]},
      {stage092[41]},
      {stage093[40], stage093[41], stage093[42], stage093[43], stage093[44], stage093[45]},
      {stage095[58], stage094[57], stage093[72], stage092[64], stage091[78]}
   );
   gpc615_5 gpc615_5_1936(
      {stage091[64], stage091[65], stage091[66], stage091[67], stage091[68]},
      {stage092[42]},
      {stage093[46], stage093[47], stage093[48], stage093[49], stage093[50], stage093[51]},
      {stage095[59], stage094[58], stage093[73], stage092[65], stage091[79]}
   );
   gpc1_1 gpc1_1_1937(
      {stage092[43]},
      {stage092[66]}
   );
   gpc1_1 gpc1_1_1938(
      {stage092[44]},
      {stage092[67]}
   );
   gpc1_1 gpc1_1_1939(
      {stage092[45]},
      {stage092[68]}
   );
   gpc1_1 gpc1_1_1940(
      {stage092[46]},
      {stage092[69]}
   );
   gpc1_1 gpc1_1_1941(
      {stage092[47]},
      {stage092[70]}
   );
   gpc1_1 gpc1_1_1942(
      {stage092[48]},
      {stage092[71]}
   );
   gpc1_1 gpc1_1_1943(
      {stage092[49]},
      {stage092[72]}
   );
   gpc1_1 gpc1_1_1944(
      {stage092[50]},
      {stage092[73]}
   );
   gpc1_1 gpc1_1_1945(
      {stage092[51]},
      {stage092[74]}
   );
   gpc1_1 gpc1_1_1946(
      {stage092[52]},
      {stage092[75]}
   );
   gpc1_1 gpc1_1_1947(
      {stage092[53]},
      {stage092[76]}
   );
   gpc1_1 gpc1_1_1948(
      {stage092[54]},
      {stage092[77]}
   );
   gpc1_1 gpc1_1_1949(
      {stage092[55]},
      {stage092[78]}
   );
   gpc1_1 gpc1_1_1950(
      {stage092[56]},
      {stage092[79]}
   );
   gpc1_1 gpc1_1_1951(
      {stage092[57]},
      {stage092[80]}
   );
   gpc1_1 gpc1_1_1952(
      {stage092[58]},
      {stage092[81]}
   );
   gpc1_1 gpc1_1_1953(
      {stage092[59]},
      {stage092[82]}
   );
   gpc1_1 gpc1_1_1954(
      {stage093[52]},
      {stage093[74]}
   );
   gpc1_1 gpc1_1_1955(
      {stage093[53]},
      {stage093[75]}
   );
   gpc1_1 gpc1_1_1956(
      {stage093[54]},
      {stage093[76]}
   );
   gpc1_1 gpc1_1_1957(
      {stage093[55]},
      {stage093[77]}
   );
   gpc1_1 gpc1_1_1958(
      {stage093[56]},
      {stage093[78]}
   );
   gpc1_1 gpc1_1_1959(
      {stage093[57]},
      {stage093[79]}
   );
   gpc615_5 gpc615_5_1960(
      {stage093[58], stage093[59], stage093[60], stage093[61], stage093[62]},
      {stage094[33]},
      {stage095[32], stage095[33], stage095[34], stage095[35], stage095[36], stage095[37]},
      {stage097[43], stage096[45], stage095[60], stage094[59], stage093[80]}
   );
   gpc615_5 gpc615_5_1961(
      {stage093[63], stage093[64], stage093[65], stage093[66], stage093[67]},
      {stage094[34]},
      {stage095[38], stage095[39], stage095[40], stage095[41], stage095[42], stage095[43]},
      {stage097[44], stage096[46], stage095[61], stage094[60], stage093[81]}
   );
   gpc1_1 gpc1_1_1962(
      {stage094[35]},
      {stage094[61]}
   );
   gpc1_1 gpc1_1_1963(
      {stage094[36]},
      {stage094[62]}
   );
   gpc1_1 gpc1_1_1964(
      {stage094[37]},
      {stage094[63]}
   );
   gpc1_1 gpc1_1_1965(
      {stage094[38]},
      {stage094[64]}
   );
   gpc1_1 gpc1_1_1966(
      {stage094[39]},
      {stage094[65]}
   );
   gpc1_1 gpc1_1_1967(
      {stage094[40]},
      {stage094[66]}
   );
   gpc1_1 gpc1_1_1968(
      {stage094[41]},
      {stage094[67]}
   );
   gpc1_1 gpc1_1_1969(
      {stage094[42]},
      {stage094[68]}
   );
   gpc1_1 gpc1_1_1970(
      {stage094[43]},
      {stage094[69]}
   );
   gpc1_1 gpc1_1_1971(
      {stage094[44]},
      {stage094[70]}
   );
   gpc615_5 gpc615_5_1972(
      {stage094[45], stage094[46], stage094[47], stage094[48], stage094[49]},
      {stage095[44]},
      {stage096[31], stage096[32], stage096[33], stage096[34], stage096[35], stage096[36]},
      {stage098[47], stage097[45], stage096[47], stage095[62], stage094[71]}
   );
   gpc615_5 gpc615_5_1973(
      {stage094[50], stage094[51], stage094[52], stage094[53], stage094[54]},
      {stage095[45]},
      {stage096[37], stage096[38], stage096[39], stage096[40], stage096[41], stage096[42]},
      {stage098[48], stage097[46], stage096[48], stage095[63], stage094[72]}
   );
   gpc1_1 gpc1_1_1974(
      {stage095[46]},
      {stage095[64]}
   );
   gpc1_1 gpc1_1_1975(
      {stage095[47]},
      {stage095[65]}
   );
   gpc1_1 gpc1_1_1976(
      {stage095[48]},
      {stage095[66]}
   );
   gpc1_1 gpc1_1_1977(
      {stage095[49]},
      {stage095[67]}
   );
   gpc1_1 gpc1_1_1978(
      {stage095[50]},
      {stage095[68]}
   );
   gpc1_1 gpc1_1_1979(
      {stage095[51]},
      {stage095[69]}
   );
   gpc1_1 gpc1_1_1980(
      {stage095[52]},
      {stage095[70]}
   );
   gpc1_1 gpc1_1_1981(
      {stage095[53]},
      {stage095[71]}
   );
   gpc1_1 gpc1_1_1982(
      {stage095[54]},
      {stage095[72]}
   );
   gpc1_1 gpc1_1_1983(
      {stage095[55]},
      {stage095[73]}
   );
   gpc1_1 gpc1_1_1984(
      {stage095[56]},
      {stage095[74]}
   );
   gpc1_1 gpc1_1_1985(
      {stage096[43]},
      {stage096[49]}
   );
   gpc1_1 gpc1_1_1986(
      {stage096[44]},
      {stage096[50]}
   );
   gpc1_1 gpc1_1_1987(
      {stage097[30]},
      {stage097[47]}
   );
   gpc1_1 gpc1_1_1988(
      {stage097[31]},
      {stage097[48]}
   );
   gpc1_1 gpc1_1_1989(
      {stage097[32]},
      {stage097[49]}
   );
   gpc1_1 gpc1_1_1990(
      {stage097[33]},
      {stage097[50]}
   );
   gpc1_1 gpc1_1_1991(
      {stage097[34]},
      {stage097[51]}
   );
   gpc1_1 gpc1_1_1992(
      {stage097[35]},
      {stage097[52]}
   );
   gpc1_1 gpc1_1_1993(
      {stage097[36]},
      {stage097[53]}
   );
   gpc1_1 gpc1_1_1994(
      {stage097[37]},
      {stage097[54]}
   );
   gpc1_1 gpc1_1_1995(
      {stage097[38]},
      {stage097[55]}
   );
   gpc1_1 gpc1_1_1996(
      {stage097[39]},
      {stage097[56]}
   );
   gpc1_1 gpc1_1_1997(
      {stage097[40]},
      {stage097[57]}
   );
   gpc1_1 gpc1_1_1998(
      {stage097[41]},
      {stage097[58]}
   );
   gpc1_1 gpc1_1_1999(
      {stage097[42]},
      {stage097[59]}
   );
   gpc1_1 gpc1_1_2000(
      {stage098[29]},
      {stage098[49]}
   );
   gpc1_1 gpc1_1_2001(
      {stage098[30]},
      {stage098[50]}
   );
   gpc1_1 gpc1_1_2002(
      {stage098[31]},
      {stage098[51]}
   );
   gpc1_1 gpc1_1_2003(
      {stage098[32]},
      {stage098[52]}
   );
   gpc1_1 gpc1_1_2004(
      {stage098[33]},
      {stage098[53]}
   );
   gpc1_1 gpc1_1_2005(
      {stage098[34]},
      {stage098[54]}
   );
   gpc606_5 gpc606_5_2006(
      {stage098[35], stage098[36], stage098[37], stage098[38], stage098[39], stage098[40]},
      {stage100[27], stage100[28], stage100[29], stage100[30], stage100[31], stage100[32]},
      {stage102[41], stage101[39], stage100[45], stage099[40], stage098[55]}
   );
   gpc606_5 gpc606_5_2007(
      {stage098[41], stage098[42], stage098[43], stage098[44], stage098[45], stage098[46]},
      {stage100[33], stage100[34], stage100[35], stage100[36], stage100[37], stage100[38]},
      {stage102[42], stage101[40], stage100[46], stage099[41], stage098[56]}
   );
   gpc606_5 gpc606_5_2008(
      {stage099[28], stage099[29], stage099[30], stage099[31], stage099[32], stage099[33]},
      {stage101[26], stage101[27], stage101[28], stage101[29], stage101[30], stage101[31]},
      {stage103[35], stage102[43], stage101[41], stage100[47], stage099[42]}
   );
   gpc606_5 gpc606_5_2009(
      {stage099[34], stage099[35], stage099[36], stage099[37], stage099[38], stage099[39]},
      {stage101[32], stage101[33], stage101[34], stage101[35], stage101[36], stage101[37]},
      {stage103[36], stage102[44], stage101[42], stage100[48], stage099[43]}
   );
   gpc1_1 gpc1_1_2010(
      {stage100[39]},
      {stage100[49]}
   );
   gpc1_1 gpc1_1_2011(
      {stage100[40]},
      {stage100[50]}
   );
   gpc1_1 gpc1_1_2012(
      {stage100[41]},
      {stage100[51]}
   );
   gpc1_1 gpc1_1_2013(
      {stage100[42]},
      {stage100[52]}
   );
   gpc1_1 gpc1_1_2014(
      {stage100[43]},
      {stage100[53]}
   );
   gpc1_1 gpc1_1_2015(
      {stage100[44]},
      {stage100[54]}
   );
   gpc1_1 gpc1_1_2016(
      {stage101[38]},
      {stage101[43]}
   );
   gpc1_1 gpc1_1_2017(
      {stage102[25]},
      {stage102[45]}
   );
   gpc1_1 gpc1_1_2018(
      {stage102[26]},
      {stage102[46]}
   );
   gpc1_1 gpc1_1_2019(
      {stage102[27]},
      {stage102[47]}
   );
   gpc1_1 gpc1_1_2020(
      {stage102[28]},
      {stage102[48]}
   );
   gpc1_1 gpc1_1_2021(
      {stage102[29]},
      {stage102[49]}
   );
   gpc1_1 gpc1_1_2022(
      {stage102[30]},
      {stage102[50]}
   );
   gpc1_1 gpc1_1_2023(
      {stage102[31]},
      {stage102[51]}
   );
   gpc1_1 gpc1_1_2024(
      {stage102[32]},
      {stage102[52]}
   );
   gpc1_1 gpc1_1_2025(
      {stage102[33]},
      {stage102[53]}
   );
   gpc1_1 gpc1_1_2026(
      {stage102[34]},
      {stage102[54]}
   );
   gpc606_5 gpc606_5_2027(
      {stage102[35], stage102[36], stage102[37], stage102[38], stage102[39], stage102[40]},
      {stage104[23], stage104[24], stage104[25], stage104[26], stage104[27], stage104[28]},
      {stage106[34], stage105[49], stage104[32], stage103[37], stage102[55]}
   );
   gpc1_1 gpc1_1_2028(
      {stage103[24]},
      {stage103[38]}
   );
   gpc1_1 gpc1_1_2029(
      {stage103[25]},
      {stage103[39]}
   );
   gpc1_1 gpc1_1_2030(
      {stage103[26]},
      {stage103[40]}
   );
   gpc1_1 gpc1_1_2031(
      {stage103[27]},
      {stage103[41]}
   );
   gpc1_1 gpc1_1_2032(
      {stage103[28]},
      {stage103[42]}
   );
   gpc1_1 gpc1_1_2033(
      {stage103[29]},
      {stage103[43]}
   );
   gpc1_1 gpc1_1_2034(
      {stage103[30]},
      {stage103[44]}
   );
   gpc1_1 gpc1_1_2035(
      {stage103[31]},
      {stage103[45]}
   );
   gpc1_1 gpc1_1_2036(
      {stage103[32]},
      {stage103[46]}
   );
   gpc1_1 gpc1_1_2037(
      {stage103[33]},
      {stage103[47]}
   );
   gpc1_1 gpc1_1_2038(
      {stage103[34]},
      {stage103[48]}
   );
   gpc1343_5 gpc1343_5_2039(
      {stage104[29], stage104[30], stage104[31]},
      {stage105[22], stage105[23], stage105[24], stage105[25]},
      {stage106[21], stage106[22], stage106[23]},
      {stage107[20]},
      {stage108[33], stage107[27], stage106[35], stage105[50], stage104[33]}
   );
   gpc1_1 gpc1_1_2040(
      {stage105[26]},
      {stage105[51]}
   );
   gpc1_1 gpc1_1_2041(
      {stage105[27]},
      {stage105[52]}
   );
   gpc1_1 gpc1_1_2042(
      {stage105[28]},
      {stage105[53]}
   );
   gpc1_1 gpc1_1_2043(
      {stage105[29]},
      {stage105[54]}
   );
   gpc1_1 gpc1_1_2044(
      {stage105[30]},
      {stage105[55]}
   );
   gpc1_1 gpc1_1_2045(
      {stage105[31]},
      {stage105[56]}
   );
   gpc1_1 gpc1_1_2046(
      {stage105[32]},
      {stage105[57]}
   );
   gpc1_1 gpc1_1_2047(
      {stage105[33]},
      {stage105[58]}
   );
   gpc1_1 gpc1_1_2048(
      {stage105[34]},
      {stage105[59]}
   );
   gpc1_1 gpc1_1_2049(
      {stage105[35]},
      {stage105[60]}
   );
   gpc1_1 gpc1_1_2050(
      {stage105[36]},
      {stage105[61]}
   );
   gpc1_1 gpc1_1_2051(
      {stage105[37]},
      {stage105[62]}
   );
   gpc1_1 gpc1_1_2052(
      {stage105[38]},
      {stage105[63]}
   );
   gpc1_1 gpc1_1_2053(
      {stage105[39]},
      {stage105[64]}
   );
   gpc1_1 gpc1_1_2054(
      {stage105[40]},
      {stage105[65]}
   );
   gpc1_1 gpc1_1_2055(
      {stage105[41]},
      {stage105[66]}
   );
   gpc1_1 gpc1_1_2056(
      {stage105[42]},
      {stage105[67]}
   );
   gpc606_5 gpc606_5_2057(
      {stage105[43], stage105[44], stage105[45], stage105[46], stage105[47], stage105[48]},
      {stage107[21], stage107[22], stage107[23], stage107[24], stage107[25], stage107[26]},
      {stage109[23], stage108[34], stage107[28], stage106[36], stage105[68]}
   );
   gpc1_1 gpc1_1_2058(
      {stage106[24]},
      {stage106[37]}
   );
   gpc1_1 gpc1_1_2059(
      {stage106[25]},
      {stage106[38]}
   );
   gpc1_1 gpc1_1_2060(
      {stage106[26]},
      {stage106[39]}
   );
   gpc1_1 gpc1_1_2061(
      {stage106[27]},
      {stage106[40]}
   );
   gpc1_1 gpc1_1_2062(
      {stage106[28]},
      {stage106[41]}
   );
   gpc1_1 gpc1_1_2063(
      {stage106[29]},
      {stage106[42]}
   );
   gpc1_1 gpc1_1_2064(
      {stage106[30]},
      {stage106[43]}
   );
   gpc1_1 gpc1_1_2065(
      {stage106[31]},
      {stage106[44]}
   );
   gpc1_1 gpc1_1_2066(
      {stage106[32]},
      {stage106[45]}
   );
   gpc1_1 gpc1_1_2067(
      {stage106[33]},
      {stage106[46]}
   );
   gpc1_1 gpc1_1_2068(
      {stage108[19]},
      {stage108[35]}
   );
   gpc1_1 gpc1_1_2069(
      {stage108[20]},
      {stage108[36]}
   );
   gpc1_1 gpc1_1_2070(
      {stage108[21]},
      {stage108[37]}
   );
   gpc1_1 gpc1_1_2071(
      {stage108[22]},
      {stage108[38]}
   );
   gpc1_1 gpc1_1_2072(
      {stage108[23]},
      {stage108[39]}
   );
   gpc1_1 gpc1_1_2073(
      {stage108[24]},
      {stage108[40]}
   );
   gpc1_1 gpc1_1_2074(
      {stage108[25]},
      {stage108[41]}
   );
   gpc1_1 gpc1_1_2075(
      {stage108[26]},
      {stage108[42]}
   );
   gpc1_1 gpc1_1_2076(
      {stage108[27]},
      {stage108[43]}
   );
   gpc1415_5 gpc1415_5_2077(
      {stage108[28], stage108[29], stage108[30], stage108[31], stage108[32]},
      {stage109[18]},
      {stage110[17], stage110[18], stage110[19], stage110[20]},
      {stage111[16]},
      {stage112[23], stage111[32], stage110[27], stage109[24], stage108[44]}
   );
   gpc1_1 gpc1_1_2078(
      {stage109[19]},
      {stage109[25]}
   );
   gpc623_5 gpc623_5_2079(
      {stage109[20], stage109[21], stage109[22]},
      {stage110[21], stage110[22]},
      {stage111[17], stage111[18], stage111[19], stage111[20], stage111[21], stage111[22]},
      {stage113[25], stage112[24], stage111[33], stage110[28], stage109[26]}
   );
   gpc615_5 gpc615_5_2080(
      {stage110[23], stage110[24], stage110[25], stage110[26], 1'h0},
      {stage111[23]},
      {stage112[15], stage112[16], stage112[17], stage112[18], stage112[19], stage112[20]},
      {stage114[17], stage113[26], stage112[25], stage111[34], stage110[29]}
   );
   gpc1_1 gpc1_1_2081(
      {stage111[24]},
      {stage111[35]}
   );
   gpc1_1 gpc1_1_2082(
      {stage111[25]},
      {stage111[36]}
   );
   gpc1_1 gpc1_1_2083(
      {stage111[26]},
      {stage111[37]}
   );
   gpc1_1 gpc1_1_2084(
      {stage111[27]},
      {stage111[38]}
   );
   gpc1_1 gpc1_1_2085(
      {stage111[28]},
      {stage111[39]}
   );
   gpc1_1 gpc1_1_2086(
      {stage111[29]},
      {stage111[40]}
   );
   gpc1_1 gpc1_1_2087(
      {stage111[30]},
      {stage111[41]}
   );
   gpc1_1 gpc1_1_2088(
      {stage111[31]},
      {stage111[42]}
   );
   gpc1_1 gpc1_1_2089(
      {stage112[21]},
      {stage112[26]}
   );
   gpc1_1 gpc1_1_2090(
      {stage112[22]},
      {stage112[27]}
   );
   gpc1_1 gpc1_1_2091(
      {stage113[14]},
      {stage113[27]}
   );
   gpc1_1 gpc1_1_2092(
      {stage113[15]},
      {stage113[28]}
   );
   gpc1_1 gpc1_1_2093(
      {stage113[16]},
      {stage113[29]}
   );
   gpc1_1 gpc1_1_2094(
      {stage113[17]},
      {stage113[30]}
   );
   gpc1_1 gpc1_1_2095(
      {stage113[18]},
      {stage113[31]}
   );
   gpc1_1 gpc1_1_2096(
      {stage113[19]},
      {stage113[32]}
   );
   gpc1_1 gpc1_1_2097(
      {stage113[20]},
      {stage113[33]}
   );
   gpc1_1 gpc1_1_2098(
      {stage113[21]},
      {stage113[34]}
   );
   gpc1_1 gpc1_1_2099(
      {stage113[22]},
      {stage113[35]}
   );
   gpc1_1 gpc1_1_2100(
      {stage113[23]},
      {stage113[36]}
   );
   gpc1_1 gpc1_1_2101(
      {stage113[24]},
      {stage113[37]}
   );
   gpc1_1 gpc1_1_2102(
      {stage114[13]},
      {stage114[18]}
   );
   gpc1_1 gpc1_1_2103(
      {stage114[14]},
      {stage114[19]}
   );
   gpc1_1 gpc1_1_2104(
      {stage114[15]},
      {stage114[20]}
   );
   gpc1_1 gpc1_1_2105(
      {stage114[16]},
      {stage114[21]}
   );
   gpc1_1 gpc1_1_2106(
      {stage115[12]},
      {stage115[27]}
   );
   gpc1_1 gpc1_1_2107(
      {stage115[13]},
      {stage115[28]}
   );
   gpc1_1 gpc1_1_2108(
      {stage115[14]},
      {stage115[29]}
   );
   gpc1_1 gpc1_1_2109(
      {stage115[15]},
      {stage115[30]}
   );
   gpc1_1 gpc1_1_2110(
      {stage115[16]},
      {stage115[31]}
   );
   gpc1_1 gpc1_1_2111(
      {stage115[17]},
      {stage115[32]}
   );
   gpc1_1 gpc1_1_2112(
      {stage115[18]},
      {stage115[33]}
   );
   gpc1_1 gpc1_1_2113(
      {stage115[19]},
      {stage115[34]}
   );
   gpc1_1 gpc1_1_2114(
      {stage115[20]},
      {stage115[35]}
   );
   gpc606_5 gpc606_5_2115(
      {stage115[21], stage115[22], stage115[23], stage115[24], stage115[25], stage115[26]},
      {stage117[10], stage117[11], stage117[12], stage117[13], stage117[14], stage117[15]},
      {stage119[17], stage118[13], stage117[20], stage116[24], stage115[36]}
   );
   gpc1_1 gpc1_1_2116(
      {stage116[11]},
      {stage116[25]}
   );
   gpc1_1 gpc1_1_2117(
      {stage116[12]},
      {stage116[26]}
   );
   gpc1_1 gpc1_1_2118(
      {stage116[13]},
      {stage116[27]}
   );
   gpc1_1 gpc1_1_2119(
      {stage116[14]},
      {stage116[28]}
   );
   gpc1_1 gpc1_1_2120(
      {stage116[15]},
      {stage116[29]}
   );
   gpc1_1 gpc1_1_2121(
      {stage116[16]},
      {stage116[30]}
   );
   gpc1_1 gpc1_1_2122(
      {stage116[17]},
      {stage116[31]}
   );
   gpc606_5 gpc606_5_2123(
      {stage116[18], stage116[19], stage116[20], stage116[21], stage116[22], stage116[23]},
      {stage118[9], stage118[10], stage118[11], stage118[12], 1'h0, 1'h0},
      {stage120[9], stage119[18], stage118[14], stage117[21], stage116[32]}
   );
   gpc606_5 gpc606_5_2124(
      {stage117[16], stage117[17], stage117[18], stage117[19], 1'h0, 1'h0},
      {stage119[8], stage119[9], stage119[10], stage119[11], stage119[12], stage119[13]},
      {stage121[11], stage120[10], stage119[19], stage118[15], stage117[22]}
   );
   gpc1_1 gpc1_1_2125(
      {stage119[14]},
      {stage119[20]}
   );
   gpc1_1 gpc1_1_2126(
      {stage119[15]},
      {stage119[21]}
   );
   gpc1_1 gpc1_1_2127(
      {stage119[16]},
      {stage119[22]}
   );
   gpc1_1 gpc1_1_2128(
      {stage120[7]},
      {stage120[11]}
   );
   gpc1_1 gpc1_1_2129(
      {stage120[8]},
      {stage120[12]}
   );
   gpc1_1 gpc1_1_2130(
      {stage121[6]},
      {stage121[12]}
   );
   gpc1_1 gpc1_1_2131(
      {stage121[7]},
      {stage121[13]}
   );
   gpc1_1 gpc1_1_2132(
      {stage121[8]},
      {stage121[14]}
   );
   gpc1_1 gpc1_1_2133(
      {stage121[9]},
      {stage121[15]}
   );
   gpc1_1 gpc1_1_2134(
      {stage121[10]},
      {stage121[16]}
   );
   gpc1_1 gpc1_1_2135(
      {stage122[5]},
      {stage122[8]}
   );
   gpc1_1 gpc1_1_2136(
      {stage122[6]},
      {stage122[9]}
   );
   gpc1_1 gpc1_1_2137(
      {stage122[7]},
      {stage122[10]}
   );
   gpc1_1 gpc1_1_2138(
      {stage123[4]},
      {stage123[6]}
   );
   gpc1_1 gpc1_1_2139(
      {stage123[5]},
      {stage123[7]}
   );
   gpc1_1 gpc1_1_2140(
      {stage124[3]},
      {stage124[6]}
   );
   gpc1_1 gpc1_1_2141(
      {stage124[4]},
      {stage124[7]}
   );
   gpc1_1 gpc1_1_2142(
      {stage124[5]},
      {stage124[8]}
   );
   gpc1_1 gpc1_1_2143(
      {stage125[2]},
      {stage125[5]}
   );
   gpc1_1 gpc1_1_2144(
      {stage125[3]},
      {stage125[6]}
   );
   gpc1_1 gpc1_1_2145(
      {stage125[4]},
      {stage125[7]}
   );
   gpc1_1 gpc1_1_2146(
      {stage126[1]},
      {stage126[2]}
   );
   gpc1_1 gpc1_1_2147(
      {stage000[2]},
      {stage000[3]}
   );
   gpc1_1 gpc1_1_2148(
      {stage001[3]},
      {stage001[4]}
   );
   gpc1_1 gpc1_1_2149(
      {stage002[4]},
      {stage002[5]}
   );
   gpc1_1 gpc1_1_2150(
      {stage003[6]},
      {stage003[8]}
   );
   gpc1_1 gpc1_1_2151(
      {stage003[7]},
      {stage003[9]}
   );
   gpc1_1 gpc1_1_2152(
      {stage004[10]},
      {stage004[11]}
   );
   gpc1_1 gpc1_1_2153(
      {stage005[13]},
      {stage005[20]}
   );
   gpc1_1 gpc1_1_2154(
      {stage005[14]},
      {stage005[21]}
   );
   gpc1_1 gpc1_1_2155(
      {stage005[15]},
      {stage005[22]}
   );
   gpc1_1 gpc1_1_2156(
      {stage005[16]},
      {stage005[23]}
   );
   gpc1_1 gpc1_1_2157(
      {stage005[17]},
      {stage005[24]}
   );
   gpc1_1 gpc1_1_2158(
      {stage005[18]},
      {stage005[25]}
   );
   gpc1_1 gpc1_1_2159(
      {stage005[19]},
      {stage005[26]}
   );
   gpc615_5 gpc615_5_2160(
      {stage006[14], stage006[15], 1'h0, 1'h0, 1'h0},
      {stage007[16]},
      {stage008[14], stage008[15], stage008[16], stage008[17], stage008[18], stage008[19]},
      {stage010[15], stage009[30], stage008[20], stage007[25], stage006[16]}
   );
   gpc1_1 gpc1_1_2161(
      {stage007[17]},
      {stage007[26]}
   );
   gpc1_1 gpc1_1_2162(
      {stage007[18]},
      {stage007[27]}
   );
   gpc606_5 gpc606_5_2163(
      {stage007[19], stage007[20], stage007[21], stage007[22], stage007[23], stage007[24]},
      {stage009[20], stage009[21], stage009[22], stage009[23], stage009[24], stage009[25]},
      {stage011[28], stage010[16], stage009[31], stage008[21], stage007[28]}
   );
   gpc1_1 gpc1_1_2164(
      {stage009[26]},
      {stage009[32]}
   );
   gpc1_1 gpc1_1_2165(
      {stage009[27]},
      {stage009[33]}
   );
   gpc1_1 gpc1_1_2166(
      {stage009[28]},
      {stage009[34]}
   );
   gpc1_1 gpc1_1_2167(
      {stage009[29]},
      {stage009[35]}
   );
   gpc1_1 gpc1_1_2168(
      {stage010[13]},
      {stage010[17]}
   );
   gpc1_1 gpc1_1_2169(
      {stage010[14]},
      {stage010[18]}
   );
   gpc1_1 gpc1_1_2170(
      {stage011[25]},
      {stage011[29]}
   );
   gpc1_1 gpc1_1_2171(
      {stage011[26]},
      {stage011[30]}
   );
   gpc1_1 gpc1_1_2172(
      {stage011[27]},
      {stage011[31]}
   );
   gpc606_5 gpc606_5_2173(
      {stage012[17], stage012[18], stage012[19], stage012[20], stage012[21], stage012[22]},
      {stage014[21], stage014[22], stage014[23], stage014[24], stage014[25], stage014[26]},
      {stage016[31], stage015[33], stage014[30], stage013[29], stage012[23]}
   );
   gpc1_1 gpc1_1_2174(
      {stage013[26]},
      {stage013[30]}
   );
   gpc1_1 gpc1_1_2175(
      {stage013[27]},
      {stage013[31]}
   );
   gpc1_1 gpc1_1_2176(
      {stage013[28]},
      {stage013[32]}
   );
   gpc1_1 gpc1_1_2177(
      {stage014[27]},
      {stage014[31]}
   );
   gpc1_1 gpc1_1_2178(
      {stage014[28]},
      {stage014[32]}
   );
   gpc1_1 gpc1_1_2179(
      {stage014[29]},
      {stage014[33]}
   );
   gpc1_1 gpc1_1_2180(
      {stage015[26]},
      {stage015[34]}
   );
   gpc606_5 gpc606_5_2181(
      {stage015[27], stage015[28], stage015[29], stage015[30], stage015[31], stage015[32]},
      {stage017[34], stage017[35], stage017[36], stage017[37], stage017[38], stage017[39]},
      {stage019[48], stage018[28], stage017[52], stage016[32], stage015[35]}
   );
   gpc1_1 gpc1_1_2182(
      {stage016[26]},
      {stage016[33]}
   );
   gpc1_1 gpc1_1_2183(
      {stage016[27]},
      {stage016[34]}
   );
   gpc1_1 gpc1_1_2184(
      {stage016[28]},
      {stage016[35]}
   );
   gpc1_1 gpc1_1_2185(
      {stage016[29]},
      {stage016[36]}
   );
   gpc1_1 gpc1_1_2186(
      {stage016[30]},
      {stage016[37]}
   );
   gpc1_1 gpc1_1_2187(
      {stage017[40]},
      {stage017[53]}
   );
   gpc1_1 gpc1_1_2188(
      {stage017[41]},
      {stage017[54]}
   );
   gpc615_5 gpc615_5_2189(
      {stage017[42], stage017[43], stage017[44], stage017[45], stage017[46]},
      {stage018[25]},
      {stage019[34], stage019[35], stage019[36], stage019[37], stage019[38], stage019[39]},
      {stage021[42], stage020[46], stage019[49], stage018[29], stage017[55]}
   );
   gpc615_5 gpc615_5_2190(
      {stage017[47], stage017[48], stage017[49], stage017[50], stage017[51]},
      {stage018[26]},
      {stage019[40], stage019[41], stage019[42], stage019[43], stage019[44], stage019[45]},
      {stage021[43], stage020[47], stage019[50], stage018[30], stage017[56]}
   );
   gpc1_1 gpc1_1_2191(
      {stage018[27]},
      {stage018[31]}
   );
   gpc1_1 gpc1_1_2192(
      {stage019[46]},
      {stage019[51]}
   );
   gpc1_1 gpc1_1_2193(
      {stage019[47]},
      {stage019[52]}
   );
   gpc606_5 gpc606_5_2194(
      {stage020[35], stage020[36], stage020[37], stage020[38], stage020[39], stage020[40]},
      {stage022[42], stage022[43], stage022[44], stage022[45], stage022[46], stage022[47]},
      {stage024[37], stage023[57], stage022[56], stage021[44], stage020[48]}
   );
   gpc615_5 gpc615_5_2195(
      {stage020[41], stage020[42], stage020[43], stage020[44], stage020[45]},
      {stage021[32]},
      {stage022[48], stage022[49], stage022[50], stage022[51], stage022[52], stage022[53]},
      {stage024[38], stage023[58], stage022[57], stage021[45], stage020[49]}
   );
   gpc623_5 gpc623_5_2196(
      {stage021[33], stage021[34], stage021[35]},
      {stage022[54], stage022[55]},
      {stage023[45], stage023[46], stage023[47], stage023[48], stage023[49], stage023[50]},
      {stage025[61], stage024[39], stage023[59], stage022[58], stage021[46]}
   );
   gpc606_5 gpc606_5_2197(
      {stage021[36], stage021[37], stage021[38], stage021[39], stage021[40], stage021[41]},
      {stage023[51], stage023[52], stage023[53], stage023[54], stage023[55], stage023[56]},
      {stage025[62], stage024[40], stage023[60], stage022[59], stage021[47]}
   );
   gpc606_5 gpc606_5_2198(
      {stage024[32], stage024[33], stage024[34], stage024[35], stage024[36], 1'h0},
      {stage026[43], stage026[44], stage026[45], stage026[46], stage026[47], stage026[48]},
      {stage028[49], stage027[79], stage026[56], stage025[63], stage024[41]}
   );
   gpc1_1 gpc1_1_2199(
      {stage025[48]},
      {stage025[64]}
   );
   gpc606_5 gpc606_5_2200(
      {stage025[49], stage025[50], stage025[51], stage025[52], stage025[53], stage025[54]},
      {stage027[52], stage027[53], stage027[54], stage027[55], stage027[56], stage027[57]},
      {stage029[61], stage028[50], stage027[80], stage026[57], stage025[65]}
   );
   gpc606_5 gpc606_5_2201(
      {stage025[55], stage025[56], stage025[57], stage025[58], stage025[59], stage025[60]},
      {stage027[58], stage027[59], stage027[60], stage027[61], stage027[62], stage027[63]},
      {stage029[62], stage028[51], stage027[81], stage026[58], stage025[66]}
   );
   gpc1_1 gpc1_1_2202(
      {stage026[49]},
      {stage026[59]}
   );
   gpc1_1 gpc1_1_2203(
      {stage026[50]},
      {stage026[60]}
   );
   gpc615_5 gpc615_5_2204(
      {stage026[51], stage026[52], stage026[53], stage026[54], stage026[55]},
      {stage027[64]},
      {stage028[41], stage028[42], stage028[43], stage028[44], stage028[45], stage028[46]},
      {stage030[56], stage029[63], stage028[52], stage027[82], stage026[61]}
   );
   gpc1_1 gpc1_1_2205(
      {stage027[65]},
      {stage027[83]}
   );
   gpc1_1 gpc1_1_2206(
      {stage027[66]},
      {stage027[84]}
   );
   gpc1_1 gpc1_1_2207(
      {stage027[67]},
      {stage027[85]}
   );
   gpc1_1 gpc1_1_2208(
      {stage027[68]},
      {stage027[86]}
   );
   gpc615_5 gpc615_5_2209(
      {stage027[69], stage027[70], stage027[71], stage027[72], stage027[73]},
      {stage028[47]},
      {stage029[49], stage029[50], stage029[51], stage029[52], stage029[53], stage029[54]},
      {stage031[59], stage030[57], stage029[64], stage028[53], stage027[87]}
   );
   gpc615_5 gpc615_5_2210(
      {stage027[74], stage027[75], stage027[76], stage027[77], stage027[78]},
      {stage028[48]},
      {stage029[55], stage029[56], stage029[57], stage029[58], stage029[59], stage029[60]},
      {stage031[60], stage030[58], stage029[65], stage028[54], stage027[88]}
   );
   gpc615_5 gpc615_5_2211(
      {stage030[46], stage030[47], stage030[48], stage030[49], stage030[50]},
      {stage031[50]},
      {stage032[66], stage032[67], stage032[68], stage032[69], stage032[70], stage032[71]},
      {stage034[66], stage033[50], stage032[87], stage031[61], stage030[59]}
   );
   gpc615_5 gpc615_5_2212(
      {stage030[51], stage030[52], stage030[53], stage030[54], stage030[55]},
      {stage031[51]},
      {stage032[72], stage032[73], stage032[74], stage032[75], stage032[76], stage032[77]},
      {stage034[67], stage033[51], stage032[88], stage031[62], stage030[60]}
   );
   gpc1_1 gpc1_1_2213(
      {stage031[52]},
      {stage031[63]}
   );
   gpc606_5 gpc606_5_2214(
      {stage031[53], stage031[54], stage031[55], stage031[56], stage031[57], stage031[58]},
      {stage033[43], stage033[44], stage033[45], stage033[46], stage033[47], stage033[48]},
      {stage035[57], stage034[68], stage033[52], stage032[89], stage031[64]}
   );
   gpc1_1 gpc1_1_2215(
      {stage032[78]},
      {stage032[90]}
   );
   gpc1_1 gpc1_1_2216(
      {stage032[79]},
      {stage032[91]}
   );
   gpc1_1 gpc1_1_2217(
      {stage032[80]},
      {stage032[92]}
   );
   gpc606_5 gpc606_5_2218(
      {stage032[81], stage032[82], stage032[83], stage032[84], stage032[85], stage032[86]},
      {stage034[58], stage034[59], stage034[60], stage034[61], stage034[62], stage034[63]},
      {stage036[61], stage035[58], stage034[69], stage033[53], stage032[93]}
   );
   gpc1_1 gpc1_1_2219(
      {stage033[49]},
      {stage033[54]}
   );
   gpc1_1 gpc1_1_2220(
      {stage034[64]},
      {stage034[70]}
   );
   gpc1_1 gpc1_1_2221(
      {stage034[65]},
      {stage034[71]}
   );
   gpc1_1 gpc1_1_2222(
      {stage035[50]},
      {stage035[59]}
   );
   gpc1_1 gpc1_1_2223(
      {stage035[51]},
      {stage035[60]}
   );
   gpc1_1 gpc1_1_2224(
      {stage035[52]},
      {stage035[61]}
   );
   gpc1_1 gpc1_1_2225(
      {stage035[53]},
      {stage035[62]}
   );
   gpc1_1 gpc1_1_2226(
      {stage035[54]},
      {stage035[63]}
   );
   gpc1_1 gpc1_1_2227(
      {stage035[55]},
      {stage035[64]}
   );
   gpc1_1 gpc1_1_2228(
      {stage035[56]},
      {stage035[65]}
   );
   gpc1_1 gpc1_1_2229(
      {stage036[49]},
      {stage036[62]}
   );
   gpc1_1 gpc1_1_2230(
      {stage036[50]},
      {stage036[63]}
   );
   gpc1_1 gpc1_1_2231(
      {stage036[51]},
      {stage036[64]}
   );
   gpc623_5 gpc623_5_2232(
      {stage036[52], stage036[53], stage036[54]},
      {stage037[55], stage037[56]},
      {stage038[64], stage038[65], stage038[66], stage038[67], stage038[68], stage038[69]},
      {stage040[74], stage039[60], stage038[84], stage037[67], stage036[65]}
   );
   gpc623_5 gpc623_5_2233(
      {stage036[55], stage036[56], stage036[57]},
      {stage037[57], stage037[58]},
      {stage038[70], stage038[71], stage038[72], stage038[73], stage038[74], stage038[75]},
      {stage040[75], stage039[61], stage038[85], stage037[68], stage036[66]}
   );
   gpc1343_5 gpc1343_5_2234(
      {stage036[58], stage036[59], stage036[60]},
      {stage037[59], stage037[60], stage037[61], stage037[62]},
      {stage038[76], stage038[77], stage038[78]},
      {stage039[56]},
      {stage040[76], stage039[62], stage038[86], stage037[69], stage036[67]}
   );
   gpc207_4 gpc207_4_2235(
      {stage037[63], stage037[64], stage037[65], stage037[66], 1'h0, 1'h0, 1'h0},
      {stage039[57], stage039[58]},
      {stage040[77], stage039[63], stage038[87], stage037[70]}
   );
   gpc606_5 gpc606_5_2236(
      {stage038[79], stage038[80], stage038[81], stage038[82], stage038[83], 1'h0},
      {stage040[56], stage040[57], stage040[58], stage040[59], stage040[60], stage040[61]},
      {stage042[79], stage041[77], stage040[78], stage039[64], stage038[88]}
   );
   gpc1_1 gpc1_1_2237(
      {stage039[59]},
      {stage039[65]}
   );
   gpc1_1 gpc1_1_2238(
      {stage040[62]},
      {stage040[79]}
   );
   gpc1_1 gpc1_1_2239(
      {stage040[63]},
      {stage040[80]}
   );
   gpc1_1 gpc1_1_2240(
      {stage040[64]},
      {stage040[81]}
   );
   gpc1_1 gpc1_1_2241(
      {stage040[65]},
      {stage040[82]}
   );
   gpc1_1 gpc1_1_2242(
      {stage040[66]},
      {stage040[83]}
   );
   gpc1_1 gpc1_1_2243(
      {stage040[67]},
      {stage040[84]}
   );
   gpc606_5 gpc606_5_2244(
      {stage040[68], stage040[69], stage040[70], stage040[71], stage040[72], stage040[73]},
      {stage042[67], stage042[68], stage042[69], stage042[70], stage042[71], stage042[72]},
      {stage044[79], stage043[83], stage042[80], stage041[78], stage040[85]}
   );
   gpc1_1 gpc1_1_2245(
      {stage041[63]},
      {stage041[79]}
   );
   gpc1_1 gpc1_1_2246(
      {stage041[64]},
      {stage041[80]}
   );
   gpc606_5 gpc606_5_2247(
      {stage041[65], stage041[66], stage041[67], stage041[68], stage041[69], stage041[70]},
      {stage043[64], stage043[65], stage043[66], stage043[67], stage043[68], stage043[69]},
      {stage045[78], stage044[80], stage043[84], stage042[81], stage041[81]}
   );
   gpc606_5 gpc606_5_2248(
      {stage041[71], stage041[72], stage041[73], stage041[74], stage041[75], stage041[76]},
      {stage043[70], stage043[71], stage043[72], stage043[73], stage043[74], stage043[75]},
      {stage045[79], stage044[81], stage043[85], stage042[82], stage041[82]}
   );
   gpc1_1 gpc1_1_2249(
      {stage042[73]},
      {stage042[83]}
   );
   gpc1_1 gpc1_1_2250(
      {stage042[74]},
      {stage042[84]}
   );
   gpc1_1 gpc1_1_2251(
      {stage042[75]},
      {stage042[85]}
   );
   gpc1_1 gpc1_1_2252(
      {stage042[76]},
      {stage042[86]}
   );
   gpc1_1 gpc1_1_2253(
      {stage042[77]},
      {stage042[87]}
   );
   gpc1_1 gpc1_1_2254(
      {stage042[78]},
      {stage042[88]}
   );
   gpc1_1 gpc1_1_2255(
      {stage043[76]},
      {stage043[86]}
   );
   gpc1_1 gpc1_1_2256(
      {stage043[77]},
      {stage043[87]}
   );
   gpc615_5 gpc615_5_2257(
      {stage043[78], stage043[79], stage043[80], stage043[81], stage043[82]},
      {stage044[72]},
      {stage045[69], stage045[70], stage045[71], stage045[72], stage045[73], stage045[74]},
      {stage047[102], stage046[82], stage045[80], stage044[82], stage043[88]}
   );
   gpc1_1 gpc1_1_2258(
      {stage044[73]},
      {stage044[83]}
   );
   gpc615_5 gpc615_5_2259(
      {stage044[74], stage044[75], stage044[76], stage044[77], stage044[78]},
      {stage045[75]},
      {stage046[64], stage046[65], stage046[66], stage046[67], stage046[68], stage046[69]},
      {stage048[118], stage047[103], stage046[83], stage045[81], stage044[84]}
   );
   gpc1_1 gpc1_1_2260(
      {stage045[76]},
      {stage045[82]}
   );
   gpc1_1 gpc1_1_2261(
      {stage045[77]},
      {stage045[83]}
   );
   gpc606_5 gpc606_5_2262(
      {stage046[70], stage046[71], stage046[72], stage046[73], stage046[74], stage046[75]},
      {stage048[87], stage048[88], stage048[89], stage048[90], stage048[91], stage048[92]},
      {stage050[89], stage049[86], stage048[119], stage047[104], stage046[84]}
   );
   gpc606_5 gpc606_5_2263(
      {stage046[76], stage046[77], stage046[78], stage046[79], stage046[80], stage046[81]},
      {stage048[93], stage048[94], stage048[95], stage048[96], stage048[97], stage048[98]},
      {stage050[90], stage049[87], stage048[120], stage047[105], stage046[85]}
   );
   gpc615_5 gpc615_5_2264(
      {stage047[92], stage047[93], stage047[94], stage047[95], stage047[96]},
      {stage048[99]},
      {stage049[72], stage049[73], stage049[74], stage049[75], stage049[76], stage049[77]},
      {stage051[78], stage050[91], stage049[88], stage048[121], stage047[106]}
   );
   gpc615_5 gpc615_5_2265(
      {stage047[97], stage047[98], stage047[99], stage047[100], stage047[101]},
      {stage048[100]},
      {stage049[78], stage049[79], stage049[80], stage049[81], stage049[82], stage049[83]},
      {stage051[79], stage050[92], stage049[89], stage048[122], stage047[107]}
   );
   gpc1_1 gpc1_1_2266(
      {stage048[101]},
      {stage048[123]}
   );
   gpc1_1 gpc1_1_2267(
      {stage048[102]},
      {stage048[124]}
   );
   gpc1_1 gpc1_1_2268(
      {stage048[103]},
      {stage048[125]}
   );
   gpc1_1 gpc1_1_2269(
      {stage048[104]},
      {stage048[126]}
   );
   gpc1_1 gpc1_1_2270(
      {stage048[105]},
      {stage048[127]}
   );
   gpc606_5 gpc606_5_2271(
      {stage048[106], stage048[107], stage048[108], stage048[109], stage048[110], stage048[111]},
      {stage050[76], stage050[77], stage050[78], stage050[79], stage050[80], stage050[81]},
      {stage052[98], stage051[80], stage050[93], stage049[90], stage048[128]}
   );
   gpc606_5 gpc606_5_2272(
      {stage048[112], stage048[113], stage048[114], stage048[115], stage048[116], stage048[117]},
      {stage050[82], stage050[83], stage050[84], stage050[85], stage050[86], stage050[87]},
      {stage052[99], stage051[81], stage050[94], stage049[91], stage048[129]}
   );
   gpc1_1 gpc1_1_2273(
      {stage049[84]},
      {stage049[92]}
   );
   gpc1_1 gpc1_1_2274(
      {stage049[85]},
      {stage049[93]}
   );
   gpc1_1 gpc1_1_2275(
      {stage050[88]},
      {stage050[95]}
   );
   gpc615_5 gpc615_5_2276(
      {stage051[68], stage051[69], stage051[70], stage051[71], stage051[72]},
      {stage052[84]},
      {stage053[101], stage053[102], stage053[103], stage053[104], stage053[105], stage053[106]},
      {stage055[104], stage054[116], stage053[123], stage052[100], stage051[82]}
   );
   gpc615_5 gpc615_5_2277(
      {stage051[73], stage051[74], stage051[75], stage051[76], stage051[77]},
      {stage052[85]},
      {stage053[107], stage053[108], stage053[109], stage053[110], stage053[111], stage053[112]},
      {stage055[105], stage054[117], stage053[124], stage052[101], stage051[83]}
   );
   gpc606_5 gpc606_5_2278(
      {stage052[86], stage052[87], stage052[88], stage052[89], stage052[90], stage052[91]},
      {stage054[100], stage054[101], stage054[102], stage054[103], stage054[104], stage054[105]},
      {stage056[87], stage055[106], stage054[118], stage053[125], stage052[102]}
   );
   gpc606_5 gpc606_5_2279(
      {stage052[92], stage052[93], stage052[94], stage052[95], stage052[96], stage052[97]},
      {stage054[106], stage054[107], stage054[108], stage054[109], stage054[110], stage054[111]},
      {stage056[88], stage055[107], stage054[119], stage053[126], stage052[103]}
   );
   gpc1_1 gpc1_1_2280(
      {stage053[113]},
      {stage053[127]}
   );
   gpc1_1 gpc1_1_2281(
      {stage053[114]},
      {stage053[128]}
   );
   gpc1_1 gpc1_1_2282(
      {stage053[115]},
      {stage053[129]}
   );
   gpc1_1 gpc1_1_2283(
      {stage053[116]},
      {stage053[130]}
   );
   gpc606_5 gpc606_5_2284(
      {stage053[117], stage053[118], stage053[119], stage053[120], stage053[121], stage053[122]},
      {stage055[84], stage055[85], stage055[86], stage055[87], stage055[88], stage055[89]},
      {stage057[89], stage056[89], stage055[108], stage054[120], stage053[131]}
   );
   gpc1_1 gpc1_1_2285(
      {stage054[112]},
      {stage054[121]}
   );
   gpc1_1 gpc1_1_2286(
      {stage054[113]},
      {stage054[122]}
   );
   gpc1_1 gpc1_1_2287(
      {stage054[114]},
      {stage054[123]}
   );
   gpc1_1 gpc1_1_2288(
      {stage054[115]},
      {stage054[124]}
   );
   gpc1_1 gpc1_1_2289(
      {stage055[90]},
      {stage055[109]}
   );
   gpc1_1 gpc1_1_2290(
      {stage055[91]},
      {stage055[110]}
   );
   gpc1_1 gpc1_1_2291(
      {stage055[92]},
      {stage055[111]}
   );
   gpc1_1 gpc1_1_2292(
      {stage055[93]},
      {stage055[112]}
   );
   gpc1_1 gpc1_1_2293(
      {stage055[94]},
      {stage055[113]}
   );
   gpc1_1 gpc1_1_2294(
      {stage055[95]},
      {stage055[114]}
   );
   gpc1_1 gpc1_1_2295(
      {stage055[96]},
      {stage055[115]}
   );
   gpc1_1 gpc1_1_2296(
      {stage055[97]},
      {stage055[116]}
   );
   gpc606_5 gpc606_5_2297(
      {stage055[98], stage055[99], stage055[100], stage055[101], stage055[102], stage055[103]},
      {stage057[79], stage057[80], stage057[81], stage057[82], stage057[83], stage057[84]},
      {stage059[103], stage058[95], stage057[90], stage056[90], stage055[117]}
   );
   gpc1_1 gpc1_1_2298(
      {stage056[75]},
      {stage056[91]}
   );
   gpc1_1 gpc1_1_2299(
      {stage056[76]},
      {stage056[92]}
   );
   gpc615_5 gpc615_5_2300(
      {stage056[77], stage056[78], stage056[79], stage056[80], stage056[81]},
      {stage057[85]},
      {stage058[83], stage058[84], stage058[85], stage058[86], stage058[87], stage058[88]},
      {stage060[99], stage059[104], stage058[96], stage057[91], stage056[93]}
   );
   gpc615_5 gpc615_5_2301(
      {stage056[82], stage056[83], stage056[84], stage056[85], stage056[86]},
      {stage057[86]},
      {stage058[89], stage058[90], stage058[91], stage058[92], stage058[93], stage058[94]},
      {stage060[100], stage059[105], stage058[97], stage057[92], stage056[94]}
   );
   gpc1_1 gpc1_1_2302(
      {stage057[87]},
      {stage057[93]}
   );
   gpc1_1 gpc1_1_2303(
      {stage057[88]},
      {stage057[94]}
   );
   gpc1_1 gpc1_1_2304(
      {stage059[91]},
      {stage059[106]}
   );
   gpc1_1 gpc1_1_2305(
      {stage059[92]},
      {stage059[107]}
   );
   gpc1_1 gpc1_1_2306(
      {stage059[93]},
      {stage059[108]}
   );
   gpc1_1 gpc1_1_2307(
      {stage059[94]},
      {stage059[109]}
   );
   gpc1_1 gpc1_1_2308(
      {stage059[95]},
      {stage059[110]}
   );
   gpc7_3 gpc7_3_2309(
      {stage059[96], stage059[97], stage059[98], stage059[99], stage059[100], stage059[101], stage059[102]},
      {stage061[120], stage060[101], stage059[111]}
   );
   gpc615_5 gpc615_5_2310(
      {stage060[85], stage060[86], stage060[87], stage060[88], stage060[89]},
      {stage061[103]},
      {stage062[102], stage062[103], stage062[104], stage062[105], stage062[106], stage062[107]},
      {stage064[108], stage063[129], stage062[126], stage061[121], stage060[102]}
   );
   gpc615_5 gpc615_5_2311(
      {stage060[90], stage060[91], stage060[92], stage060[93], stage060[94]},
      {stage061[104]},
      {stage062[108], stage062[109], stage062[110], stage062[111], stage062[112], stage062[113]},
      {stage064[109], stage063[130], stage062[127], stage061[122], stage060[103]}
   );
   gpc615_5 gpc615_5_2312(
      {stage060[95], stage060[96], stage060[97], stage060[98], 1'h0},
      {stage061[105]},
      {stage062[114], stage062[115], stage062[116], stage062[117], stage062[118], stage062[119]},
      {stage064[110], stage063[131], stage062[128], stage061[123], stage060[104]}
   );
   gpc1_1 gpc1_1_2313(
      {stage061[106]},
      {stage061[124]}
   );
   gpc1_1 gpc1_1_2314(
      {stage061[107]},
      {stage061[125]}
   );
   gpc1_1 gpc1_1_2315(
      {stage061[108]},
      {stage061[126]}
   );
   gpc1_1 gpc1_1_2316(
      {stage061[109]},
      {stage061[127]}
   );
   gpc615_5 gpc615_5_2317(
      {stage061[110], stage061[111], stage061[112], stage061[113], stage061[114]},
      {stage062[120]},
      {stage063[104], stage063[105], stage063[106], stage063[107], stage063[108], stage063[109]},
      {stage065[116], stage064[111], stage063[132], stage062[129], stage061[128]}
   );
   gpc615_5 gpc615_5_2318(
      {stage061[115], stage061[116], stage061[117], stage061[118], stage061[119]},
      {stage062[121]},
      {stage063[110], stage063[111], stage063[112], stage063[113], stage063[114], stage063[115]},
      {stage065[117], stage064[112], stage063[133], stage062[130], stage061[129]}
   );
   gpc1_1 gpc1_1_2319(
      {stage062[122]},
      {stage062[131]}
   );
   gpc1_1 gpc1_1_2320(
      {stage062[123]},
      {stage062[132]}
   );
   gpc1_1 gpc1_1_2321(
      {stage062[124]},
      {stage062[133]}
   );
   gpc1_1 gpc1_1_2322(
      {stage062[125]},
      {stage062[134]}
   );
   gpc1_1 gpc1_1_2323(
      {stage063[116]},
      {stage063[134]}
   );
   gpc1_1 gpc1_1_2324(
      {stage063[117]},
      {stage063[135]}
   );
   gpc606_5 gpc606_5_2325(
      {stage063[118], stage063[119], stage063[120], stage063[121], stage063[122], stage063[123]},
      {stage065[91], stage065[92], stage065[93], stage065[94], stage065[95], stage065[96]},
      {stage067[115], stage066[99], stage065[118], stage064[113], stage063[136]}
   );
   gpc615_5 gpc615_5_2326(
      {stage063[124], stage063[125], stage063[126], stage063[127], stage063[128]},
      {stage064[97]},
      {stage065[97], stage065[98], stage065[99], stage065[100], stage065[101], stage065[102]},
      {stage067[116], stage066[100], stage065[119], stage064[114], stage063[137]}
   );
   gpc615_5 gpc615_5_2327(
      {stage064[98], stage064[99], stage064[100], stage064[101], stage064[102]},
      {stage065[103]},
      {stage066[85], stage066[86], stage066[87], stage066[88], stage066[89], stage066[90]},
      {stage068[99], stage067[117], stage066[101], stage065[120], stage064[115]}
   );
   gpc615_5 gpc615_5_2328(
      {stage064[103], stage064[104], stage064[105], stage064[106], stage064[107]},
      {stage065[104]},
      {stage066[91], stage066[92], stage066[93], stage066[94], stage066[95], stage066[96]},
      {stage068[100], stage067[118], stage066[102], stage065[121], stage064[116]}
   );
   gpc606_5 gpc606_5_2329(
      {stage065[105], stage065[106], stage065[107], stage065[108], stage065[109], stage065[110]},
      {stage067[103], stage067[104], stage067[105], stage067[106], stage067[107], stage067[108]},
      {stage069[107], stage068[101], stage067[119], stage066[103], stage065[122]}
   );
   gpc615_5 gpc615_5_2330(
      {stage065[111], stage065[112], stage065[113], stage065[114], stage065[115]},
      {stage066[97]},
      {stage067[109], stage067[110], stage067[111], stage067[112], stage067[113], stage067[114]},
      {stage069[108], stage068[102], stage067[120], stage066[104], stage065[123]}
   );
   gpc1_1 gpc1_1_2331(
      {stage066[98]},
      {stage066[105]}
   );
   gpc1_1 gpc1_1_2332(
      {stage068[85]},
      {stage068[103]}
   );
   gpc1_1 gpc1_1_2333(
      {stage068[86]},
      {stage068[104]}
   );
   gpc615_5 gpc615_5_2334(
      {stage068[87], stage068[88], stage068[89], stage068[90], stage068[91]},
      {stage069[92]},
      {stage070[90], stage070[91], stage070[92], stage070[93], stage070[94], stage070[95]},
      {stage072[99], stage071[100], stage070[102], stage069[109], stage068[105]}
   );
   gpc207_4 gpc207_4_2335(
      {stage068[92], stage068[93], stage068[94], stage068[95], stage068[96], stage068[97], stage068[98]},
      {stage070[96], stage070[97]},
      {stage071[101], stage070[103], stage069[110], stage068[106]}
   );
   gpc1_1 gpc1_1_2336(
      {stage069[93]},
      {stage069[111]}
   );
   gpc1_1 gpc1_1_2337(
      {stage069[94]},
      {stage069[112]}
   );
   gpc1_1 gpc1_1_2338(
      {stage069[95]},
      {stage069[113]}
   );
   gpc1_1 gpc1_1_2339(
      {stage069[96]},
      {stage069[114]}
   );
   gpc615_5 gpc615_5_2340(
      {stage069[97], stage069[98], stage069[99], stage069[100], stage069[101]},
      {stage070[98]},
      {stage071[80], stage071[81], stage071[82], stage071[83], stage071[84], stage071[85]},
      {stage073[92], stage072[100], stage071[102], stage070[104], stage069[115]}
   );
   gpc615_5 gpc615_5_2341(
      {stage069[102], stage069[103], stage069[104], stage069[105], stage069[106]},
      {stage070[99]},
      {stage071[86], stage071[87], stage071[88], stage071[89], stage071[90], stage071[91]},
      {stage073[93], stage072[101], stage071[103], stage070[105], stage069[116]}
   );
   gpc1_1 gpc1_1_2342(
      {stage070[100]},
      {stage070[106]}
   );
   gpc1_1 gpc1_1_2343(
      {stage070[101]},
      {stage070[107]}
   );
   gpc1_1 gpc1_1_2344(
      {stage071[92]},
      {stage071[104]}
   );
   gpc1_1 gpc1_1_2345(
      {stage071[93]},
      {stage071[105]}
   );
   gpc1_1 gpc1_1_2346(
      {stage071[94]},
      {stage071[106]}
   );
   gpc1_1 gpc1_1_2347(
      {stage071[95]},
      {stage071[107]}
   );
   gpc1_1 gpc1_1_2348(
      {stage071[96]},
      {stage071[108]}
   );
   gpc1_1 gpc1_1_2349(
      {stage071[97]},
      {stage071[109]}
   );
   gpc1_1 gpc1_1_2350(
      {stage071[98]},
      {stage071[110]}
   );
   gpc1_1 gpc1_1_2351(
      {stage071[99]},
      {stage071[111]}
   );
   gpc1_1 gpc1_1_2352(
      {stage072[83]},
      {stage072[102]}
   );
   gpc615_5 gpc615_5_2353(
      {stage072[84], stage072[85], stage072[86], stage072[87], stage072[88]},
      {stage073[84]},
      {stage074[81], stage074[82], stage074[83], stage074[84], stage074[85], stage074[86]},
      {stage076[84], stage075[88], stage074[105], stage073[94], stage072[103]}
   );
   gpc615_5 gpc615_5_2354(
      {stage072[89], stage072[90], stage072[91], stage072[92], stage072[93]},
      {stage073[85]},
      {stage074[87], stage074[88], stage074[89], stage074[90], stage074[91], stage074[92]},
      {stage076[85], stage075[89], stage074[106], stage073[95], stage072[104]}
   );
   gpc615_5 gpc615_5_2355(
      {stage072[94], stage072[95], stage072[96], stage072[97], stage072[98]},
      {stage073[86]},
      {stage074[93], stage074[94], stage074[95], stage074[96], stage074[97], stage074[98]},
      {stage076[86], stage075[90], stage074[107], stage073[96], stage072[105]}
   );
   gpc615_5 gpc615_5_2356(
      {stage073[87], stage073[88], stage073[89], stage073[90], stage073[91]},
      {stage074[99]},
      {stage075[78], stage075[79], stage075[80], stage075[81], stage075[82], stage075[83]},
      {stage077[90], stage076[87], stage075[91], stage074[108], stage073[97]}
   );
   gpc1_1 gpc1_1_2357(
      {stage074[100]},
      {stage074[109]}
   );
   gpc1_1 gpc1_1_2358(
      {stage074[101]},
      {stage074[110]}
   );
   gpc1_1 gpc1_1_2359(
      {stage074[102]},
      {stage074[111]}
   );
   gpc1_1 gpc1_1_2360(
      {stage074[103]},
      {stage074[112]}
   );
   gpc1_1 gpc1_1_2361(
      {stage074[104]},
      {stage074[113]}
   );
   gpc1_1 gpc1_1_2362(
      {stage075[84]},
      {stage075[92]}
   );
   gpc1_1 gpc1_1_2363(
      {stage075[85]},
      {stage075[93]}
   );
   gpc1_1 gpc1_1_2364(
      {stage075[86]},
      {stage075[94]}
   );
   gpc1_1 gpc1_1_2365(
      {stage075[87]},
      {stage075[95]}
   );
   gpc1_1 gpc1_1_2366(
      {stage076[73]},
      {stage076[88]}
   );
   gpc615_5 gpc615_5_2367(
      {stage076[74], stage076[75], stage076[76], stage076[77], stage076[78]},
      {stage077[75]},
      {stage078[71], stage078[72], stage078[73], stage078[74], stage078[75], stage078[76]},
      {stage080[85], stage079[101], stage078[89], stage077[91], stage076[89]}
   );
   gpc615_5 gpc615_5_2368(
      {stage076[79], stage076[80], stage076[81], stage076[82], stage076[83]},
      {stage077[76]},
      {stage078[77], stage078[78], stage078[79], stage078[80], stage078[81], stage078[82]},
      {stage080[86], stage079[102], stage078[90], stage077[92], stage076[90]}
   );
   gpc1_1 gpc1_1_2369(
      {stage077[77]},
      {stage077[93]}
   );
   gpc1_1 gpc1_1_2370(
      {stage077[78]},
      {stage077[94]}
   );
   gpc1_1 gpc1_1_2371(
      {stage077[79]},
      {stage077[95]}
   );
   gpc615_5 gpc615_5_2372(
      {stage077[80], stage077[81], stage077[82], stage077[83], stage077[84]},
      {stage078[83]},
      {stage079[85], stage079[86], stage079[87], stage079[88], stage079[89], stage079[90]},
      {stage081[84], stage080[87], stage079[103], stage078[91], stage077[96]}
   );
   gpc2135_5 gpc2135_5_2373(
      {stage077[85], stage077[86], stage077[87], stage077[88], stage077[89]},
      {stage078[84], stage078[85], stage078[86]},
      {stage079[91]},
      {stage080[71], stage080[72]},
      {stage081[85], stage080[88], stage079[104], stage078[92], stage077[97]}
   );
   gpc1_1 gpc1_1_2374(
      {stage078[87]},
      {stage078[93]}
   );
   gpc1_1 gpc1_1_2375(
      {stage078[88]},
      {stage078[94]}
   );
   gpc1_1 gpc1_1_2376(
      {stage079[92]},
      {stage079[105]}
   );
   gpc1_1 gpc1_1_2377(
      {stage079[93]},
      {stage079[106]}
   );
   gpc1_1 gpc1_1_2378(
      {stage079[94]},
      {stage079[107]}
   );
   gpc1_1 gpc1_1_2379(
      {stage079[95]},
      {stage079[108]}
   );
   gpc1_1 gpc1_1_2380(
      {stage079[96]},
      {stage079[109]}
   );
   gpc1_1 gpc1_1_2381(
      {stage079[97]},
      {stage079[110]}
   );
   gpc1_1 gpc1_1_2382(
      {stage079[98]},
      {stage079[111]}
   );
   gpc1_1 gpc1_1_2383(
      {stage079[99]},
      {stage079[112]}
   );
   gpc1_1 gpc1_1_2384(
      {stage079[100]},
      {stage079[113]}
   );
   gpc1_1 gpc1_1_2385(
      {stage080[73]},
      {stage080[89]}
   );
   gpc1_1 gpc1_1_2386(
      {stage080[74]},
      {stage080[90]}
   );
   gpc615_5 gpc615_5_2387(
      {stage080[75], stage080[76], stage080[77], stage080[78], stage080[79]},
      {stage081[75]},
      {stage082[66], stage082[67], stage082[68], stage082[69], stage082[70], stage082[71]},
      {stage084[84], stage083[74], stage082[78], stage081[86], stage080[91]}
   );
   gpc615_5 gpc615_5_2388(
      {stage080[80], stage080[81], stage080[82], stage080[83], stage080[84]},
      {stage081[76]},
      {stage082[72], stage082[73], stage082[74], stage082[75], stage082[76], stage082[77]},
      {stage084[85], stage083[75], stage082[79], stage081[87], stage080[92]}
   );
   gpc1_1 gpc1_1_2389(
      {stage081[77]},
      {stage081[88]}
   );
   gpc1_1 gpc1_1_2390(
      {stage081[78]},
      {stage081[89]}
   );
   gpc1_1 gpc1_1_2391(
      {stage081[79]},
      {stage081[90]}
   );
   gpc1_1 gpc1_1_2392(
      {stage081[80]},
      {stage081[91]}
   );
   gpc1_1 gpc1_1_2393(
      {stage081[81]},
      {stage081[92]}
   );
   gpc1_1 gpc1_1_2394(
      {stage081[82]},
      {stage081[93]}
   );
   gpc1_1 gpc1_1_2395(
      {stage081[83]},
      {stage081[94]}
   );
   gpc1_1 gpc1_1_2396(
      {stage083[63]},
      {stage083[76]}
   );
   gpc1_1 gpc1_1_2397(
      {stage083[64]},
      {stage083[77]}
   );
   gpc1_1 gpc1_1_2398(
      {stage083[65]},
      {stage083[78]}
   );
   gpc1_1 gpc1_1_2399(
      {stage083[66]},
      {stage083[79]}
   );
   gpc7_3 gpc7_3_2400(
      {stage083[67], stage083[68], stage083[69], stage083[70], stage083[71], stage083[72], stage083[73]},
      {stage085[81], stage084[86], stage083[80]}
   );
   gpc1_1 gpc1_1_2401(
      {stage084[74]},
      {stage084[87]}
   );
   gpc1343_5 gpc1343_5_2402(
      {stage084[75], stage084[76], stage084[77]},
      {stage085[68], stage085[69], stage085[70], stage085[71]},
      {stage086[66], stage086[67], stage086[68]},
      {stage087[54]},
      {stage088[66], stage087[64], stage086[81], stage085[82], stage084[88]}
   );
   gpc1343_5 gpc1343_5_2403(
      {stage084[78], stage084[79], stage084[80]},
      {stage085[72], stage085[73], stage085[74], stage085[75]},
      {stage086[69], stage086[70], stage086[71]},
      {stage087[55]},
      {stage088[67], stage087[65], stage086[82], stage085[83], stage084[89]}
   );
   gpc1343_5 gpc1343_5_2404(
      {stage084[81], stage084[82], stage084[83]},
      {stage085[76], stage085[77], stage085[78], stage085[79]},
      {stage086[72], stage086[73], stage086[74]},
      {stage087[56]},
      {stage088[68], stage087[66], stage086[83], stage085[84], stage084[90]}
   );
   gpc1_1 gpc1_1_2405(
      {stage085[80]},
      {stage085[85]}
   );
   gpc606_5 gpc606_5_2406(
      {stage086[75], stage086[76], stage086[77], stage086[78], stage086[79], stage086[80]},
      {stage088[53], stage088[54], stage088[55], stage088[56], stage088[57], stage088[58]},
      {stage090[67], stage089[71], stage088[69], stage087[67], stage086[84]}
   );
   gpc1_1 gpc1_1_2407(
      {stage087[57]},
      {stage087[68]}
   );
   gpc1_1 gpc1_1_2408(
      {stage087[58]},
      {stage087[69]}
   );
   gpc615_5 gpc615_5_2409(
      {stage087[59], stage087[60], stage087[61], stage087[62], stage087[63]},
      {stage088[59]},
      {stage089[60], stage089[61], stage089[62], stage089[63], stage089[64], stage089[65]},
      {stage091[80], stage090[68], stage089[72], stage088[70], stage087[70]}
   );
   gpc1_1 gpc1_1_2410(
      {stage088[60]},
      {stage088[71]}
   );
   gpc615_5 gpc615_5_2411(
      {stage088[61], stage088[62], stage088[63], stage088[64], stage088[65]},
      {stage089[66]},
      {stage090[53], stage090[54], stage090[55], stage090[56], stage090[57], stage090[58]},
      {stage092[83], stage091[81], stage090[69], stage089[73], stage088[72]}
   );
   gpc1_1 gpc1_1_2412(
      {stage089[67]},
      {stage089[74]}
   );
   gpc1_1 gpc1_1_2413(
      {stage089[68]},
      {stage089[75]}
   );
   gpc1_1 gpc1_1_2414(
      {stage089[69]},
      {stage089[76]}
   );
   gpc1_1 gpc1_1_2415(
      {stage089[70]},
      {stage089[77]}
   );
   gpc1_1 gpc1_1_2416(
      {stage090[59]},
      {stage090[70]}
   );
   gpc1_1 gpc1_1_2417(
      {stage090[60]},
      {stage090[71]}
   );
   gpc1_1 gpc1_1_2418(
      {stage090[61]},
      {stage090[72]}
   );
   gpc615_5 gpc615_5_2419(
      {stage090[62], stage090[63], stage090[64], stage090[65], stage090[66]},
      {stage091[69]},
      {stage092[60], stage092[61], stage092[62], stage092[63], stage092[64], stage092[65]},
      {stage094[73], stage093[82], stage092[84], stage091[82], stage090[73]}
   );
   gpc615_5 gpc615_5_2420(
      {stage091[70], stage091[71], stage091[72], stage091[73], stage091[74]},
      {stage092[66]},
      {stage093[68], stage093[69], stage093[70], stage093[71], stage093[72], stage093[73]},
      {stage095[75], stage094[74], stage093[83], stage092[85], stage091[83]}
   );
   gpc615_5 gpc615_5_2421(
      {stage091[75], stage091[76], stage091[77], stage091[78], stage091[79]},
      {stage092[67]},
      {stage093[74], stage093[75], stage093[76], stage093[77], stage093[78], stage093[79]},
      {stage095[76], stage094[75], stage093[84], stage092[86], stage091[84]}
   );
   gpc1_1 gpc1_1_2422(
      {stage092[68]},
      {stage092[87]}
   );
   gpc1_1 gpc1_1_2423(
      {stage092[69]},
      {stage092[88]}
   );
   gpc1_1 gpc1_1_2424(
      {stage092[70]},
      {stage092[89]}
   );
   gpc606_5 gpc606_5_2425(
      {stage092[71], stage092[72], stage092[73], stage092[74], stage092[75], stage092[76]},
      {stage094[55], stage094[56], stage094[57], stage094[58], stage094[59], stage094[60]},
      {stage096[51], stage095[77], stage094[76], stage093[85], stage092[90]}
   );
   gpc606_5 gpc606_5_2426(
      {stage092[77], stage092[78], stage092[79], stage092[80], stage092[81], stage092[82]},
      {stage094[61], stage094[62], stage094[63], stage094[64], stage094[65], stage094[66]},
      {stage096[52], stage095[78], stage094[77], stage093[86], stage092[91]}
   );
   gpc1_1 gpc1_1_2427(
      {stage093[80]},
      {stage093[87]}
   );
   gpc1_1 gpc1_1_2428(
      {stage093[81]},
      {stage093[88]}
   );
   gpc606_5 gpc606_5_2429(
      {stage094[67], stage094[68], stage094[69], stage094[70], stage094[71], stage094[72]},
      {stage096[45], stage096[46], stage096[47], stage096[48], stage096[49], stage096[50]},
      {stage098[57], stage097[60], stage096[53], stage095[79], stage094[78]}
   );
   gpc606_5 gpc606_5_2430(
      {stage095[57], stage095[58], stage095[59], stage095[60], stage095[61], stage095[62]},
      {stage097[43], stage097[44], stage097[45], stage097[46], stage097[47], stage097[48]},
      {stage099[44], stage098[58], stage097[61], stage096[54], stage095[80]}
   );
   gpc606_5 gpc606_5_2431(
      {stage095[63], stage095[64], stage095[65], stage095[66], stage095[67], stage095[68]},
      {stage097[49], stage097[50], stage097[51], stage097[52], stage097[53], stage097[54]},
      {stage099[45], stage098[59], stage097[62], stage096[55], stage095[81]}
   );
   gpc606_5 gpc606_5_2432(
      {stage095[69], stage095[70], stage095[71], stage095[72], stage095[73], stage095[74]},
      {stage097[55], stage097[56], stage097[57], stage097[58], stage097[59], 1'h0},
      {stage099[46], stage098[60], stage097[63], stage096[56], stage095[82]}
   );
   gpc1_1 gpc1_1_2433(
      {stage098[47]},
      {stage098[61]}
   );
   gpc1_1 gpc1_1_2434(
      {stage098[48]},
      {stage098[62]}
   );
   gpc1_1 gpc1_1_2435(
      {stage098[49]},
      {stage098[63]}
   );
   gpc1_1 gpc1_1_2436(
      {stage098[50]},
      {stage098[64]}
   );
   gpc1_1 gpc1_1_2437(
      {stage098[51]},
      {stage098[65]}
   );
   gpc1_1 gpc1_1_2438(
      {stage098[52]},
      {stage098[66]}
   );
   gpc1_1 gpc1_1_2439(
      {stage098[53]},
      {stage098[67]}
   );
   gpc1_1 gpc1_1_2440(
      {stage098[54]},
      {stage098[68]}
   );
   gpc1_1 gpc1_1_2441(
      {stage098[55]},
      {stage098[69]}
   );
   gpc1_1 gpc1_1_2442(
      {stage098[56]},
      {stage098[70]}
   );
   gpc1_1 gpc1_1_2443(
      {stage099[40]},
      {stage099[47]}
   );
   gpc1_1 gpc1_1_2444(
      {stage099[41]},
      {stage099[48]}
   );
   gpc1_1 gpc1_1_2445(
      {stage099[42]},
      {stage099[49]}
   );
   gpc1_1 gpc1_1_2446(
      {stage099[43]},
      {stage099[50]}
   );
   gpc1_1 gpc1_1_2447(
      {stage100[45]},
      {stage100[55]}
   );
   gpc1_1 gpc1_1_2448(
      {stage100[46]},
      {stage100[56]}
   );
   gpc1_1 gpc1_1_2449(
      {stage100[47]},
      {stage100[57]}
   );
   gpc1_1 gpc1_1_2450(
      {stage100[48]},
      {stage100[58]}
   );
   gpc1_1 gpc1_1_2451(
      {stage100[49]},
      {stage100[59]}
   );
   gpc615_5 gpc615_5_2452(
      {stage100[50], stage100[51], stage100[52], stage100[53], stage100[54]},
      {stage101[39]},
      {stage102[41], stage102[42], stage102[43], stage102[44], stage102[45], stage102[46]},
      {stage104[34], stage103[49], stage102[56], stage101[44], stage100[60]}
   );
   gpc615_5 gpc615_5_2453(
      {stage101[40], stage101[41], stage101[42], stage101[43], 1'h0},
      {stage102[47]},
      {stage103[35], stage103[36], stage103[37], stage103[38], stage103[39], stage103[40]},
      {stage105[69], stage104[35], stage103[50], stage102[57], stage101[45]}
   );
   gpc1_1 gpc1_1_2454(
      {stage102[48]},
      {stage102[58]}
   );
   gpc1_1 gpc1_1_2455(
      {stage102[49]},
      {stage102[59]}
   );
   gpc1_1 gpc1_1_2456(
      {stage102[50]},
      {stage102[60]}
   );
   gpc1_1 gpc1_1_2457(
      {stage102[51]},
      {stage102[61]}
   );
   gpc1_1 gpc1_1_2458(
      {stage102[52]},
      {stage102[62]}
   );
   gpc1_1 gpc1_1_2459(
      {stage102[53]},
      {stage102[63]}
   );
   gpc1_1 gpc1_1_2460(
      {stage102[54]},
      {stage102[64]}
   );
   gpc1_1 gpc1_1_2461(
      {stage102[55]},
      {stage102[65]}
   );
   gpc615_5 gpc615_5_2462(
      {stage103[41], stage103[42], stage103[43], stage103[44], stage103[45]},
      {stage104[32]},
      {stage105[49], stage105[50], stage105[51], stage105[52], stage105[53], stage105[54]},
      {stage107[29], stage106[47], stage105[70], stage104[36], stage103[51]}
   );
   gpc615_5 gpc615_5_2463(
      {stage103[46], stage103[47], stage103[48], 1'h0, 1'h0},
      {stage104[33]},
      {stage105[55], stage105[56], stage105[57], stage105[58], stage105[59], stage105[60]},
      {stage107[30], stage106[48], stage105[71], stage104[37], stage103[52]}
   );
   gpc1_1 gpc1_1_2464(
      {stage105[61]},
      {stage105[72]}
   );
   gpc1_1 gpc1_1_2465(
      {stage105[62]},
      {stage105[73]}
   );
   gpc1_1 gpc1_1_2466(
      {stage105[63]},
      {stage105[74]}
   );
   gpc2135_5 gpc2135_5_2467(
      {stage105[64], stage105[65], stage105[66], stage105[67], stage105[68]},
      {stage106[34], stage106[35], stage106[36]},
      {stage107[27]},
      {stage108[33], stage108[34]},
      {stage109[27], stage108[45], stage107[31], stage106[49], stage105[75]}
   );
   gpc1_1 gpc1_1_2468(
      {stage106[37]},
      {stage106[50]}
   );
   gpc1_1 gpc1_1_2469(
      {stage106[38]},
      {stage106[51]}
   );
   gpc1_1 gpc1_1_2470(
      {stage106[39]},
      {stage106[52]}
   );
   gpc1_1 gpc1_1_2471(
      {stage106[40]},
      {stage106[53]}
   );
   gpc606_5 gpc606_5_2472(
      {stage106[41], stage106[42], stage106[43], stage106[44], stage106[45], stage106[46]},
      {stage108[35], stage108[36], stage108[37], stage108[38], stage108[39], stage108[40]},
      {stage110[30], stage109[28], stage108[46], stage107[32], stage106[54]}
   );
   gpc1_1 gpc1_1_2473(
      {stage107[28]},
      {stage107[33]}
   );
   gpc1_1 gpc1_1_2474(
      {stage108[41]},
      {stage108[47]}
   );
   gpc1_1 gpc1_1_2475(
      {stage108[42]},
      {stage108[48]}
   );
   gpc1_1 gpc1_1_2476(
      {stage108[43]},
      {stage108[49]}
   );
   gpc1_1 gpc1_1_2477(
      {stage108[44]},
      {stage108[50]}
   );
   gpc1_1 gpc1_1_2478(
      {stage109[23]},
      {stage109[29]}
   );
   gpc1343_5 gpc1343_5_2479(
      {stage109[24], stage109[25], stage109[26]},
      {stage110[27], stage110[28], stage110[29], 1'h0},
      {stage111[32], stage111[33], stage111[34]},
      {stage112[23]},
      {stage113[38], stage112[28], stage111[43], stage110[31], stage109[30]}
   );
   gpc615_5 gpc615_5_2480(
      {stage111[35], stage111[36], stage111[37], stage111[38], stage111[39]},
      {stage112[24]},
      {stage113[25], stage113[26], stage113[27], stage113[28], stage113[29], stage113[30]},
      {stage115[37], stage114[22], stage113[39], stage112[29], stage111[44]}
   );
   gpc1325_5 gpc1325_5_2481(
      {stage111[40], stage111[41], stage111[42], 1'h0, 1'h0},
      {stage112[25], stage112[26]},
      {stage113[31], stage113[32], stage113[33]},
      {stage114[17]},
      {stage115[38], stage114[23], stage113[40], stage112[30], stage111[45]}
   );
   gpc1_1 gpc1_1_2482(
      {stage112[27]},
      {stage112[31]}
   );
   gpc606_5 gpc606_5_2483(
      {stage113[34], stage113[35], stage113[36], stage113[37], 1'h0, 1'h0},
      {stage115[27], stage115[28], stage115[29], stage115[30], stage115[31], stage115[32]},
      {stage117[23], stage116[33], stage115[39], stage114[24], stage113[41]}
   );
   gpc1_1 gpc1_1_2484(
      {stage114[18]},
      {stage114[25]}
   );
   gpc1_1 gpc1_1_2485(
      {stage114[19]},
      {stage114[26]}
   );
   gpc1_1 gpc1_1_2486(
      {stage114[20]},
      {stage114[27]}
   );
   gpc1_1 gpc1_1_2487(
      {stage114[21]},
      {stage114[28]}
   );
   gpc1_1 gpc1_1_2488(
      {stage115[33]},
      {stage115[40]}
   );
   gpc1_1 gpc1_1_2489(
      {stage115[34]},
      {stage115[41]}
   );
   gpc1_1 gpc1_1_2490(
      {stage115[35]},
      {stage115[42]}
   );
   gpc1_1 gpc1_1_2491(
      {stage115[36]},
      {stage115[43]}
   );
   gpc1_1 gpc1_1_2492(
      {stage116[24]},
      {stage116[34]}
   );
   gpc1_1 gpc1_1_2493(
      {stage116[25]},
      {stage116[35]}
   );
   gpc1_1 gpc1_1_2494(
      {stage116[26]},
      {stage116[36]}
   );
   gpc1_1 gpc1_1_2495(
      {stage116[27]},
      {stage116[37]}
   );
   gpc1415_5 gpc1415_5_2496(
      {stage116[28], stage116[29], stage116[30], stage116[31], stage116[32]},
      {stage117[20]},
      {stage118[13], stage118[14], stage118[15], 1'h0},
      {stage119[17]},
      {stage120[13], stage119[23], stage118[16], stage117[24], stage116[38]}
   );
   gpc1_1 gpc1_1_2497(
      {stage117[21]},
      {stage117[25]}
   );
   gpc1_1 gpc1_1_2498(
      {stage117[22]},
      {stage117[26]}
   );
   gpc606_5 gpc606_5_2499(
      {stage119[18], stage119[19], stage119[20], stage119[21], stage119[22], 1'h0},
      {stage121[11], stage121[12], stage121[13], stage121[14], stage121[15], stage121[16]},
      {stage123[8], stage122[11], stage121[17], stage120[14], stage119[24]}
   );
   gpc1_1 gpc1_1_2500(
      {stage120[9]},
      {stage120[15]}
   );
   gpc1_1 gpc1_1_2501(
      {stage120[10]},
      {stage120[16]}
   );
   gpc1_1 gpc1_1_2502(
      {stage120[11]},
      {stage120[17]}
   );
   gpc1_1 gpc1_1_2503(
      {stage120[12]},
      {stage120[18]}
   );
   gpc1_1 gpc1_1_2504(
      {stage122[8]},
      {stage122[12]}
   );
   gpc1_1 gpc1_1_2505(
      {stage122[9]},
      {stage122[13]}
   );
   gpc1_1 gpc1_1_2506(
      {stage122[10]},
      {stage122[14]}
   );
   gpc1_1 gpc1_1_2507(
      {stage123[6]},
      {stage123[9]}
   );
   gpc1_1 gpc1_1_2508(
      {stage123[7]},
      {stage123[10]}
   );
   gpc1_1 gpc1_1_2509(
      {stage124[6]},
      {stage124[9]}
   );
   gpc1_1 gpc1_1_2510(
      {stage124[7]},
      {stage124[10]}
   );
   gpc1_1 gpc1_1_2511(
      {stage124[8]},
      {stage124[11]}
   );
   gpc1406_5 gpc1406_5_2512(
      {stage125[5], stage125[6], stage125[7], 1'h0, 1'h0, 1'h0},
      {1'h0, 1'h0, 1'h0, 1'h0},
      {1'h0},
      {stage128[0], stage127[0], stage126[3], stage125[8]}
   );
   gpc1_1 gpc1_1_2513(
      {stage126[2]},
      {stage126[4]}
   );
   gpc1_1 gpc1_1_2514(
      {stage000[3]},
      {stage000[4]}
   );
   gpc1_1 gpc1_1_2515(
      {stage001[4]},
      {stage001[5]}
   );
   gpc1_1 gpc1_1_2516(
      {stage002[5]},
      {stage002[6]}
   );
   gpc623_5 gpc623_5_2517(
      {stage003[8], stage003[9], 1'h0},
      {stage004[11], 1'h0},
      {stage005[20], stage005[21], stage005[22], stage005[23], stage005[24], stage005[25]},
      {stage007[29], stage006[17], stage005[27], stage004[12], stage003[10]}
   );
   gpc1_1 gpc1_1_2518(
      {stage005[26]},
      {stage005[28]}
   );
   gpc1_1 gpc1_1_2519(
      {stage006[16]},
      {stage006[18]}
   );
   gpc1_1 gpc1_1_2520(
      {stage007[25]},
      {stage007[30]}
   );
   gpc1_1 gpc1_1_2521(
      {stage007[26]},
      {stage007[31]}
   );
   gpc1_1 gpc1_1_2522(
      {stage007[27]},
      {stage007[32]}
   );
   gpc1_1 gpc1_1_2523(
      {stage007[28]},
      {stage007[33]}
   );
   gpc606_5 gpc606_5_2524(
      {stage008[20], stage008[21], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage010[15], stage010[16], stage010[17], stage010[18], 1'h0, 1'h0},
      {stage012[24], stage011[32], stage010[19], stage009[36], stage008[22]}
   );
   gpc1_1 gpc1_1_2525(
      {stage009[30]},
      {stage009[37]}
   );
   gpc1_1 gpc1_1_2526(
      {stage009[31]},
      {stage009[38]}
   );
   gpc1_1 gpc1_1_2527(
      {stage009[32]},
      {stage009[39]}
   );
   gpc1_1 gpc1_1_2528(
      {stage009[33]},
      {stage009[40]}
   );
   gpc1_1 gpc1_1_2529(
      {stage009[34]},
      {stage009[41]}
   );
   gpc1_1 gpc1_1_2530(
      {stage009[35]},
      {stage009[42]}
   );
   gpc1_1 gpc1_1_2531(
      {stage011[28]},
      {stage011[33]}
   );
   gpc1_1 gpc1_1_2532(
      {stage011[29]},
      {stage011[34]}
   );
   gpc1_1 gpc1_1_2533(
      {stage011[30]},
      {stage011[35]}
   );
   gpc1_1 gpc1_1_2534(
      {stage011[31]},
      {stage011[36]}
   );
   gpc1_1 gpc1_1_2535(
      {stage012[23]},
      {stage012[25]}
   );
   gpc1_1 gpc1_1_2536(
      {stage013[29]},
      {stage013[33]}
   );
   gpc1_1 gpc1_1_2537(
      {stage013[30]},
      {stage013[34]}
   );
   gpc1_1 gpc1_1_2538(
      {stage013[31]},
      {stage013[35]}
   );
   gpc1_1 gpc1_1_2539(
      {stage013[32]},
      {stage013[36]}
   );
   gpc606_5 gpc606_5_2540(
      {stage014[30], stage014[31], stage014[32], stage014[33], 1'h0, 1'h0},
      {stage016[31], stage016[32], stage016[33], stage016[34], stage016[35], stage016[36]},
      {stage018[32], stage017[57], stage016[38], stage015[36], stage014[34]}
   );
   gpc1_1 gpc1_1_2541(
      {stage015[33]},
      {stage015[37]}
   );
   gpc1_1 gpc1_1_2542(
      {stage015[34]},
      {stage015[38]}
   );
   gpc1_1 gpc1_1_2543(
      {stage015[35]},
      {stage015[39]}
   );
   gpc1_1 gpc1_1_2544(
      {stage016[37]},
      {stage016[39]}
   );
   gpc1_1 gpc1_1_2545(
      {stage017[52]},
      {stage017[58]}
   );
   gpc1_1 gpc1_1_2546(
      {stage017[53]},
      {stage017[59]}
   );
   gpc1_1 gpc1_1_2547(
      {stage017[54]},
      {stage017[60]}
   );
   gpc1_1 gpc1_1_2548(
      {stage017[55]},
      {stage017[61]}
   );
   gpc1_1 gpc1_1_2549(
      {stage017[56]},
      {stage017[62]}
   );
   gpc1_1 gpc1_1_2550(
      {stage018[28]},
      {stage018[33]}
   );
   gpc1_1 gpc1_1_2551(
      {stage018[29]},
      {stage018[34]}
   );
   gpc1_1 gpc1_1_2552(
      {stage018[30]},
      {stage018[35]}
   );
   gpc1_1 gpc1_1_2553(
      {stage018[31]},
      {stage018[36]}
   );
   gpc615_5 gpc615_5_2554(
      {stage019[48], stage019[49], stage019[50], stage019[51], stage019[52]},
      {stage020[46]},
      {stage021[42], stage021[43], stage021[44], stage021[45], stage021[46], stage021[47]},
      {stage023[61], stage022[60], stage021[48], stage020[50], stage019[53]}
   );
   gpc1_1 gpc1_1_2555(
      {stage020[47]},
      {stage020[51]}
   );
   gpc1_1 gpc1_1_2556(
      {stage020[48]},
      {stage020[52]}
   );
   gpc1_1 gpc1_1_2557(
      {stage020[49]},
      {stage020[53]}
   );
   gpc1_1 gpc1_1_2558(
      {stage022[56]},
      {stage022[61]}
   );
   gpc1_1 gpc1_1_2559(
      {stage022[57]},
      {stage022[62]}
   );
   gpc1_1 gpc1_1_2560(
      {stage022[58]},
      {stage022[63]}
   );
   gpc1_1 gpc1_1_2561(
      {stage022[59]},
      {stage022[64]}
   );
   gpc606_5 gpc606_5_2562(
      {stage023[57], stage023[58], stage023[59], stage023[60], 1'h0, 1'h0},
      {stage025[61], stage025[62], stage025[63], stage025[64], stage025[65], stage025[66]},
      {stage027[89], stage026[62], stage025[67], stage024[42], stage023[62]}
   );
   gpc1_1 gpc1_1_2563(
      {stage024[37]},
      {stage024[43]}
   );
   gpc1_1 gpc1_1_2564(
      {stage024[38]},
      {stage024[44]}
   );
   gpc1_1 gpc1_1_2565(
      {stage024[39]},
      {stage024[45]}
   );
   gpc1_1 gpc1_1_2566(
      {stage024[40]},
      {stage024[46]}
   );
   gpc1_1 gpc1_1_2567(
      {stage024[41]},
      {stage024[47]}
   );
   gpc606_5 gpc606_5_2568(
      {stage026[56], stage026[57], stage026[58], stage026[59], stage026[60], stage026[61]},
      {stage028[49], stage028[50], stage028[51], stage028[52], stage028[53], stage028[54]},
      {stage030[61], stage029[66], stage028[55], stage027[90], stage026[63]}
   );
   gpc1_1 gpc1_1_2569(
      {stage027[79]},
      {stage027[91]}
   );
   gpc1_1 gpc1_1_2570(
      {stage027[80]},
      {stage027[92]}
   );
   gpc1_1 gpc1_1_2571(
      {stage027[81]},
      {stage027[93]}
   );
   gpc1_1 gpc1_1_2572(
      {stage027[82]},
      {stage027[94]}
   );
   gpc606_5 gpc606_5_2573(
      {stage027[83], stage027[84], stage027[85], stage027[86], stage027[87], stage027[88]},
      {stage029[61], stage029[62], stage029[63], stage029[64], stage029[65], 1'h0},
      {stage031[65], stage030[62], stage029[67], stage028[56], stage027[95]}
   );
   gpc615_5 gpc615_5_2574(
      {stage030[56], stage030[57], stage030[58], stage030[59], stage030[60]},
      {stage031[59]},
      {stage032[87], stage032[88], stage032[89], stage032[90], stage032[91], stage032[92]},
      {stage034[72], stage033[55], stage032[94], stage031[66], stage030[63]}
   );
   gpc1_1 gpc1_1_2575(
      {stage031[60]},
      {stage031[67]}
   );
   gpc1_1 gpc1_1_2576(
      {stage031[61]},
      {stage031[68]}
   );
   gpc1_1 gpc1_1_2577(
      {stage031[62]},
      {stage031[69]}
   );
   gpc1_1 gpc1_1_2578(
      {stage031[63]},
      {stage031[70]}
   );
   gpc1_1 gpc1_1_2579(
      {stage031[64]},
      {stage031[71]}
   );
   gpc1_1 gpc1_1_2580(
      {stage032[93]},
      {stage032[95]}
   );
   gpc606_5 gpc606_5_2581(
      {stage033[50], stage033[51], stage033[52], stage033[53], stage033[54], 1'h0},
      {stage035[57], stage035[58], stage035[59], stage035[60], stage035[61], stage035[62]},
      {stage037[71], stage036[68], stage035[66], stage034[73], stage033[56]}
   );
   gpc606_5 gpc606_5_2582(
      {stage034[66], stage034[67], stage034[68], stage034[69], stage034[70], stage034[71]},
      {stage036[61], stage036[62], stage036[63], stage036[64], stage036[65], stage036[66]},
      {stage038[89], stage037[72], stage036[69], stage035[67], stage034[74]}
   );
   gpc1_1 gpc1_1_2583(
      {stage035[63]},
      {stage035[68]}
   );
   gpc1_1 gpc1_1_2584(
      {stage035[64]},
      {stage035[69]}
   );
   gpc1_1 gpc1_1_2585(
      {stage035[65]},
      {stage035[70]}
   );
   gpc1_1 gpc1_1_2586(
      {stage036[67]},
      {stage036[70]}
   );
   gpc1_1 gpc1_1_2587(
      {stage037[67]},
      {stage037[73]}
   );
   gpc1_1 gpc1_1_2588(
      {stage037[68]},
      {stage037[74]}
   );
   gpc1_1 gpc1_1_2589(
      {stage037[69]},
      {stage037[75]}
   );
   gpc1_1 gpc1_1_2590(
      {stage037[70]},
      {stage037[76]}
   );
   gpc615_5 gpc615_5_2591(
      {stage038[84], stage038[85], stage038[86], stage038[87], stage038[88]},
      {stage039[60]},
      {stage040[74], stage040[75], stage040[76], stage040[77], stage040[78], stage040[79]},
      {stage042[89], stage041[83], stage040[86], stage039[66], stage038[90]}
   );
   gpc1_1 gpc1_1_2592(
      {stage039[61]},
      {stage039[67]}
   );
   gpc1_1 gpc1_1_2593(
      {stage039[62]},
      {stage039[68]}
   );
   gpc1_1 gpc1_1_2594(
      {stage039[63]},
      {stage039[69]}
   );
   gpc1_1 gpc1_1_2595(
      {stage039[64]},
      {stage039[70]}
   );
   gpc1_1 gpc1_1_2596(
      {stage039[65]},
      {stage039[71]}
   );
   gpc1_1 gpc1_1_2597(
      {stage040[80]},
      {stage040[87]}
   );
   gpc615_5 gpc615_5_2598(
      {stage040[81], stage040[82], stage040[83], stage040[84], stage040[85]},
      {stage041[77]},
      {stage042[79], stage042[80], stage042[81], stage042[82], stage042[83], stage042[84]},
      {stage044[85], stage043[89], stage042[90], stage041[84], stage040[88]}
   );
   gpc606_5 gpc606_5_2599(
      {stage041[78], stage041[79], stage041[80], stage041[81], stage041[82], 1'h0},
      {stage043[83], stage043[84], stage043[85], stage043[86], stage043[87], stage043[88]},
      {stage045[84], stage044[86], stage043[90], stage042[91], stage041[85]}
   );
   gpc1_1 gpc1_1_2600(
      {stage042[85]},
      {stage042[92]}
   );
   gpc1_1 gpc1_1_2601(
      {stage042[86]},
      {stage042[93]}
   );
   gpc1_1 gpc1_1_2602(
      {stage042[87]},
      {stage042[94]}
   );
   gpc1_1 gpc1_1_2603(
      {stage042[88]},
      {stage042[95]}
   );
   gpc1_1 gpc1_1_2604(
      {stage044[79]},
      {stage044[87]}
   );
   gpc2135_5 gpc2135_5_2605(
      {stage044[80], stage044[81], stage044[82], stage044[83], stage044[84]},
      {stage045[78], stage045[79], stage045[80]},
      {stage046[82]},
      {stage047[102], stage047[103]},
      {stage048[130], stage047[108], stage046[86], stage045[85], stage044[88]}
   );
   gpc1_1 gpc1_1_2606(
      {stage045[81]},
      {stage045[86]}
   );
   gpc1_1 gpc1_1_2607(
      {stage045[82]},
      {stage045[87]}
   );
   gpc1_1 gpc1_1_2608(
      {stage045[83]},
      {stage045[88]}
   );
   gpc623_5 gpc623_5_2609(
      {stage046[83], stage046[84], stage046[85]},
      {stage047[104], stage047[105]},
      {stage048[118], stage048[119], stage048[120], stage048[121], stage048[122], stage048[123]},
      {stage050[96], stage049[94], stage048[131], stage047[109], stage046[87]}
   );
   gpc1_1 gpc1_1_2610(
      {stage047[106]},
      {stage047[110]}
   );
   gpc1_1 gpc1_1_2611(
      {stage047[107]},
      {stage047[111]}
   );
   gpc606_5 gpc606_5_2612(
      {stage048[124], stage048[125], stage048[126], stage048[127], stage048[128], stage048[129]},
      {stage050[89], stage050[90], stage050[91], stage050[92], stage050[93], stage050[94]},
      {stage052[104], stage051[84], stage050[97], stage049[95], stage048[132]}
   );
   gpc1_1 gpc1_1_2613(
      {stage049[86]},
      {stage049[96]}
   );
   gpc1_1 gpc1_1_2614(
      {stage049[87]},
      {stage049[97]}
   );
   gpc1_1 gpc1_1_2615(
      {stage049[88]},
      {stage049[98]}
   );
   gpc615_5 gpc615_5_2616(
      {stage049[89], stage049[90], stage049[91], stage049[92], stage049[93]},
      {stage050[95]},
      {stage051[78], stage051[79], stage051[80], stage051[81], stage051[82], stage051[83]},
      {stage053[132], stage052[105], stage051[85], stage050[98], stage049[99]}
   );
   gpc606_5 gpc606_5_2617(
      {stage052[98], stage052[99], stage052[100], stage052[101], stage052[102], stage052[103]},
      {stage054[116], stage054[117], stage054[118], stage054[119], stage054[120], stage054[121]},
      {stage056[95], stage055[118], stage054[125], stage053[133], stage052[106]}
   );
   gpc1_1 gpc1_1_2618(
      {stage053[123]},
      {stage053[134]}
   );
   gpc1_1 gpc1_1_2619(
      {stage053[124]},
      {stage053[135]}
   );
   gpc1_1 gpc1_1_2620(
      {stage053[125]},
      {stage053[136]}
   );
   gpc606_5 gpc606_5_2621(
      {stage053[126], stage053[127], stage053[128], stage053[129], stage053[130], stage053[131]},
      {stage055[104], stage055[105], stage055[106], stage055[107], stage055[108], stage055[109]},
      {stage057[95], stage056[96], stage055[119], stage054[126], stage053[137]}
   );
   gpc623_5 gpc623_5_2622(
      {stage054[122], stage054[123], stage054[124]},
      {stage055[110], stage055[111]},
      {stage056[87], stage056[88], stage056[89], stage056[90], stage056[91], stage056[92]},
      {stage058[98], stage057[96], stage056[97], stage055[120], stage054[127]}
   );
   gpc606_5 gpc606_5_2623(
      {stage055[112], stage055[113], stage055[114], stage055[115], stage055[116], stage055[117]},
      {stage057[89], stage057[90], stage057[91], stage057[92], stage057[93], stage057[94]},
      {stage059[112], stage058[99], stage057[97], stage056[98], stage055[121]}
   );
   gpc1_1 gpc1_1_2624(
      {stage056[93]},
      {stage056[99]}
   );
   gpc1_1 gpc1_1_2625(
      {stage056[94]},
      {stage056[100]}
   );
   gpc3_2 gpc3_2_2626(
      {stage058[95], stage058[96], stage058[97]},
      {stage059[113], stage058[100]}
   );
   gpc2135_5 gpc2135_5_2627(
      {stage059[103], stage059[104], stage059[105], stage059[106], stage059[107]},
      {stage060[99], stage060[100], stage060[101]},
      {stage061[120]},
      {stage062[126], stage062[127]},
      {stage063[138], stage062[135], stage061[130], stage060[105], stage059[114]}
   );
   gpc2135_5 gpc2135_5_2628(
      {stage059[108], stage059[109], stage059[110], stage059[111], 1'h0},
      {stage060[102], stage060[103], stage060[104]},
      {stage061[121]},
      {stage062[128], stage062[129]},
      {stage063[139], stage062[136], stage061[131], stage060[106], stage059[115]}
   );
   gpc1_1 gpc1_1_2629(
      {stage061[122]},
      {stage061[132]}
   );
   gpc1_1 gpc1_1_2630(
      {stage061[123]},
      {stage061[133]}
   );
   gpc606_5 gpc606_5_2631(
      {stage061[124], stage061[125], stage061[126], stage061[127], stage061[128], stage061[129]},
      {stage063[129], stage063[130], stage063[131], stage063[132], stage063[133], stage063[134]},
      {stage065[124], stage064[117], stage063[140], stage062[137], stage061[134]}
   );
   gpc615_5 gpc615_5_2632(
      {stage062[130], stage062[131], stage062[132], stage062[133], stage062[134]},
      {stage063[135]},
      {stage064[108], stage064[109], stage064[110], stage064[111], stage064[112], stage064[113]},
      {stage066[106], stage065[125], stage064[118], stage063[141], stage062[138]}
   );
   gpc1_1 gpc1_1_2633(
      {stage063[136]},
      {stage063[142]}
   );
   gpc1_1 gpc1_1_2634(
      {stage063[137]},
      {stage063[143]}
   );
   gpc623_5 gpc623_5_2635(
      {stage064[114], stage064[115], stage064[116]},
      {stage065[116], stage065[117]},
      {stage066[99], stage066[100], stage066[101], stage066[102], stage066[103], stage066[104]},
      {stage068[107], stage067[121], stage066[107], stage065[126], stage064[119]}
   );
   gpc606_5 gpc606_5_2636(
      {stage065[118], stage065[119], stage065[120], stage065[121], stage065[122], stage065[123]},
      {stage067[115], stage067[116], stage067[117], stage067[118], stage067[119], stage067[120]},
      {stage069[117], stage068[108], stage067[122], stage066[108], stage065[127]}
   );
   gpc1_1 gpc1_1_2637(
      {stage066[105]},
      {stage066[109]}
   );
   gpc1_1 gpc1_1_2638(
      {stage068[99]},
      {stage068[109]}
   );
   gpc1_1 gpc1_1_2639(
      {stage068[100]},
      {stage068[110]}
   );
   gpc1_1 gpc1_1_2640(
      {stage068[101]},
      {stage068[111]}
   );
   gpc2135_5 gpc2135_5_2641(
      {stage068[102], stage068[103], stage068[104], stage068[105], stage068[106]},
      {stage069[107], stage069[108], stage069[109]},
      {stage070[102]},
      {stage071[100], stage071[101]},
      {stage072[106], stage071[112], stage070[108], stage069[118], stage068[112]}
   );
   gpc1_1 gpc1_1_2642(
      {stage069[110]},
      {stage069[119]}
   );
   gpc1_1 gpc1_1_2643(
      {stage069[111]},
      {stage069[120]}
   );
   gpc615_5 gpc615_5_2644(
      {stage069[112], stage069[113], stage069[114], stage069[115], stage069[116]},
      {stage070[103]},
      {stage071[102], stage071[103], stage071[104], stage071[105], stage071[106], stage071[107]},
      {stage073[98], stage072[107], stage071[113], stage070[109], stage069[121]}
   );
   gpc615_5 gpc615_5_2645(
      {stage070[104], stage070[105], stage070[106], stage070[107], 1'h0},
      {stage071[108]},
      {stage072[99], stage072[100], stage072[101], stage072[102], stage072[103], stage072[104]},
      {stage074[114], stage073[99], stage072[108], stage071[114], stage070[110]}
   );
   gpc1_1 gpc1_1_2646(
      {stage071[109]},
      {stage071[115]}
   );
   gpc1_1 gpc1_1_2647(
      {stage071[110]},
      {stage071[116]}
   );
   gpc1_1 gpc1_1_2648(
      {stage071[111]},
      {stage071[117]}
   );
   gpc1_1 gpc1_1_2649(
      {stage072[105]},
      {stage072[109]}
   );
   gpc207_4 gpc207_4_2650(
      {stage073[92], stage073[93], stage073[94], stage073[95], stage073[96], stage073[97], 1'h0},
      {stage075[88], stage075[89]},
      {stage076[91], stage075[96], stage074[115], stage073[100]}
   );
   gpc1_1 gpc1_1_2651(
      {stage074[105]},
      {stage074[116]}
   );
   gpc1_1 gpc1_1_2652(
      {stage074[106]},
      {stage074[117]}
   );
   gpc1_1 gpc1_1_2653(
      {stage074[107]},
      {stage074[118]}
   );
   gpc606_5 gpc606_5_2654(
      {stage074[108], stage074[109], stage074[110], stage074[111], stage074[112], stage074[113]},
      {stage076[84], stage076[85], stage076[86], stage076[87], stage076[88], stage076[89]},
      {stage078[95], stage077[98], stage076[92], stage075[97], stage074[119]}
   );
   gpc606_5 gpc606_5_2655(
      {stage075[90], stage075[91], stage075[92], stage075[93], stage075[94], stage075[95]},
      {stage077[90], stage077[91], stage077[92], stage077[93], stage077[94], stage077[95]},
      {stage079[114], stage078[96], stage077[99], stage076[93], stage075[98]}
   );
   gpc1_1 gpc1_1_2656(
      {stage076[90]},
      {stage076[94]}
   );
   gpc1_1 gpc1_1_2657(
      {stage077[96]},
      {stage077[100]}
   );
   gpc1_1 gpc1_1_2658(
      {stage077[97]},
      {stage077[101]}
   );
   gpc1_1 gpc1_1_2659(
      {stage078[89]},
      {stage078[97]}
   );
   gpc1_1 gpc1_1_2660(
      {stage078[90]},
      {stage078[98]}
   );
   gpc1_1 gpc1_1_2661(
      {stage078[91]},
      {stage078[99]}
   );
   gpc623_5 gpc623_5_2662(
      {stage078[92], stage078[93], stage078[94]},
      {stage079[101], stage079[102]},
      {stage080[85], stage080[86], stage080[87], stage080[88], stage080[89], stage080[90]},
      {stage082[80], stage081[95], stage080[93], stage079[115], stage078[100]}
   );
   gpc1_1 gpc1_1_2663(
      {stage079[103]},
      {stage079[116]}
   );
   gpc1415_5 gpc1415_5_2664(
      {stage079[104], stage079[105], stage079[106], stage079[107], stage079[108]},
      {stage080[91]},
      {stage081[84], stage081[85], stage081[86], stage081[87]},
      {stage082[78]},
      {stage083[81], stage082[81], stage081[96], stage080[94], stage079[117]}
   );
   gpc1415_5 gpc1415_5_2665(
      {stage079[109], stage079[110], stage079[111], stage079[112], stage079[113]},
      {stage080[92]},
      {stage081[88], stage081[89], stage081[90], stage081[91]},
      {stage082[79]},
      {stage083[82], stage082[82], stage081[97], stage080[95], stage079[118]}
   );
   gpc1_1 gpc1_1_2666(
      {stage081[92]},
      {stage081[98]}
   );
   gpc1_1 gpc1_1_2667(
      {stage081[93]},
      {stage081[99]}
   );
   gpc1_1 gpc1_1_2668(
      {stage081[94]},
      {stage081[100]}
   );
   gpc1_1 gpc1_1_2669(
      {stage083[74]},
      {stage083[83]}
   );
   gpc1_1 gpc1_1_2670(
      {stage083[75]},
      {stage083[84]}
   );
   gpc1_1 gpc1_1_2671(
      {stage083[76]},
      {stage083[85]}
   );
   gpc1_1 gpc1_1_2672(
      {stage083[77]},
      {stage083[86]}
   );
   gpc623_5 gpc623_5_2673(
      {stage083[78], stage083[79], stage083[80]},
      {stage084[84], stage084[85]},
      {stage085[81], stage085[82], stage085[83], stage085[84], stage085[85], 1'h0},
      {stage087[71], stage086[85], stage085[86], stage084[91], stage083[87]}
   );
   gpc1406_5 gpc1406_5_2674(
      {stage084[86], stage084[87], stage084[88], stage084[89], stage084[90], 1'h0},
      {stage086[81], stage086[82], stage086[83], stage086[84]},
      {stage087[64]},
      {stage088[73], stage087[72], stage086[86], stage085[87], stage084[92]}
   );
   gpc223_4 gpc223_4_2675(
      {stage087[65], stage087[66], stage087[67]},
      {stage088[66], stage088[67]},
      {stage089[71], stage089[72]},
      {stage090[74], stage089[78], stage088[74], stage087[73]}
   );
   gpc223_4 gpc223_4_2676(
      {stage087[68], stage087[69], stage087[70]},
      {stage088[68], stage088[69]},
      {stage089[73], stage089[74]},
      {stage090[75], stage089[79], stage088[75], stage087[74]}
   );
   gpc623_5 gpc623_5_2677(
      {stage088[70], stage088[71], stage088[72]},
      {stage089[75], stage089[76]},
      {stage090[67], stage090[68], stage090[69], stage090[70], stage090[71], stage090[72]},
      {stage092[92], stage091[85], stage090[76], stage089[80], stage088[76]}
   );
   gpc1_1 gpc1_1_2678(
      {stage089[77]},
      {stage089[81]}
   );
   gpc1_1 gpc1_1_2679(
      {stage090[73]},
      {stage090[77]}
   );
   gpc606_5 gpc606_5_2680(
      {stage091[80], stage091[81], stage091[82], stage091[83], stage091[84], 1'h0},
      {stage093[82], stage093[83], stage093[84], stage093[85], stage093[86], stage093[87]},
      {stage095[83], stage094[79], stage093[89], stage092[93], stage091[86]}
   );
   gpc1_1 gpc1_1_2681(
      {stage092[83]},
      {stage092[94]}
   );
   gpc1_1 gpc1_1_2682(
      {stage092[84]},
      {stage092[95]}
   );
   gpc1_1 gpc1_1_2683(
      {stage092[85]},
      {stage092[96]}
   );
   gpc606_5 gpc606_5_2684(
      {stage092[86], stage092[87], stage092[88], stage092[89], stage092[90], stage092[91]},
      {stage094[73], stage094[74], stage094[75], stage094[76], stage094[77], stage094[78]},
      {stage096[57], stage095[84], stage094[80], stage093[90], stage092[97]}
   );
   gpc1_1 gpc1_1_2685(
      {stage093[88]},
      {stage093[91]}
   );
   gpc1_1 gpc1_1_2686(
      {stage095[75]},
      {stage095[85]}
   );
   gpc7_3 gpc7_3_2687(
      {stage095[76], stage095[77], stage095[78], stage095[79], stage095[80], stage095[81], stage095[82]},
      {stage097[64], stage096[58], stage095[86]}
   );
   gpc606_5 gpc606_5_2688(
      {stage096[51], stage096[52], stage096[53], stage096[54], stage096[55], stage096[56]},
      {stage098[57], stage098[58], stage098[59], stage098[60], stage098[61], stage098[62]},
      {stage100[61], stage099[51], stage098[71], stage097[65], stage096[59]}
   );
   gpc1_1 gpc1_1_2689(
      {stage097[60]},
      {stage097[66]}
   );
   gpc623_5 gpc623_5_2690(
      {stage097[61], stage097[62], stage097[63]},
      {stage098[63], stage098[64]},
      {stage099[44], stage099[45], stage099[46], stage099[47], stage099[48], stage099[49]},
      {stage101[46], stage100[62], stage099[52], stage098[72], stage097[67]}
   );
   gpc1_1 gpc1_1_2691(
      {stage098[65]},
      {stage098[73]}
   );
   gpc615_5 gpc615_5_2692(
      {stage098[66], stage098[67], stage098[68], stage098[69], stage098[70]},
      {stage099[50]},
      {stage100[55], stage100[56], stage100[57], stage100[58], stage100[59], stage100[60]},
      {stage102[66], stage101[47], stage100[63], stage099[53], stage098[74]}
   );
   gpc1_1 gpc1_1_2693(
      {stage101[44]},
      {stage101[48]}
   );
   gpc1_1 gpc1_1_2694(
      {stage101[45]},
      {stage101[49]}
   );
   gpc1_1 gpc1_1_2695(
      {stage102[56]},
      {stage102[67]}
   );
   gpc1_1 gpc1_1_2696(
      {stage102[57]},
      {stage102[68]}
   );
   gpc1_1 gpc1_1_2697(
      {stage102[58]},
      {stage102[69]}
   );
   gpc1_1 gpc1_1_2698(
      {stage102[59]},
      {stage102[70]}
   );
   gpc606_5 gpc606_5_2699(
      {stage102[60], stage102[61], stage102[62], stage102[63], stage102[64], stage102[65]},
      {stage104[34], stage104[35], stage104[36], stage104[37], 1'h0, 1'h0},
      {stage106[55], stage105[76], stage104[38], stage103[53], stage102[71]}
   );
   gpc1_1 gpc1_1_2700(
      {stage103[49]},
      {stage103[54]}
   );
   gpc1_1 gpc1_1_2701(
      {stage103[50]},
      {stage103[55]}
   );
   gpc1_1 gpc1_1_2702(
      {stage103[51]},
      {stage103[56]}
   );
   gpc1_1 gpc1_1_2703(
      {stage103[52]},
      {stage103[57]}
   );
   gpc1_1 gpc1_1_2704(
      {stage105[69]},
      {stage105[77]}
   );
   gpc1_1 gpc1_1_2705(
      {stage105[70]},
      {stage105[78]}
   );
   gpc615_5 gpc615_5_2706(
      {stage105[71], stage105[72], stage105[73], stage105[74], stage105[75]},
      {stage106[47]},
      {stage107[29], stage107[30], stage107[31], stage107[32], stage107[33], 1'h0},
      {stage109[31], stage108[51], stage107[34], stage106[56], stage105[79]}
   );
   gpc1_1 gpc1_1_2707(
      {stage106[48]},
      {stage106[57]}
   );
   gpc606_5 gpc606_5_2708(
      {stage106[49], stage106[50], stage106[51], stage106[52], stage106[53], stage106[54]},
      {stage108[45], stage108[46], stage108[47], stage108[48], stage108[49], stage108[50]},
      {stage110[32], stage109[32], stage108[52], stage107[35], stage106[58]}
   );
   gpc1_1 gpc1_1_2709(
      {stage109[27]},
      {stage109[33]}
   );
   gpc1_1 gpc1_1_2710(
      {stage109[28]},
      {stage109[34]}
   );
   gpc1_1 gpc1_1_2711(
      {stage109[29]},
      {stage109[35]}
   );
   gpc1_1 gpc1_1_2712(
      {stage109[30]},
      {stage109[36]}
   );
   gpc1_1 gpc1_1_2713(
      {stage110[30]},
      {stage110[33]}
   );
   gpc1_1 gpc1_1_2714(
      {stage110[31]},
      {stage110[34]}
   );
   gpc1343_5 gpc1343_5_2715(
      {stage111[43], stage111[44], stage111[45]},
      {stage112[28], stage112[29], stage112[30], stage112[31]},
      {stage113[38], stage113[39], stage113[40]},
      {stage114[22]},
      {stage115[44], stage114[29], stage113[42], stage112[32], stage111[46]}
   );
   gpc1_1 gpc1_1_2716(
      {stage113[41]},
      {stage113[43]}
   );
   gpc606_5 gpc606_5_2717(
      {stage114[23], stage114[24], stage114[25], stage114[26], stage114[27], stage114[28]},
      {stage116[33], stage116[34], stage116[35], stage116[36], stage116[37], stage116[38]},
      {stage118[17], stage117[27], stage116[39], stage115[45], stage114[30]}
   );
   gpc1_1 gpc1_1_2718(
      {stage115[37]},
      {stage115[46]}
   );
   gpc606_5 gpc606_5_2719(
      {stage115[38], stage115[39], stage115[40], stage115[41], stage115[42], stage115[43]},
      {stage117[23], stage117[24], stage117[25], stage117[26], 1'h0, 1'h0},
      {stage119[25], stage118[18], stage117[28], stage116[40], stage115[47]}
   );
   gpc1_1 gpc1_1_2720(
      {stage118[16]},
      {stage118[19]}
   );
   gpc1_1 gpc1_1_2721(
      {stage119[23]},
      {stage119[26]}
   );
   gpc1_1 gpc1_1_2722(
      {stage119[24]},
      {stage119[27]}
   );
   gpc606_5 gpc606_5_2723(
      {stage120[13], stage120[14], stage120[15], stage120[16], stage120[17], stage120[18]},
      {stage122[11], stage122[12], stage122[13], stage122[14], 1'h0, 1'h0},
      {stage124[12], stage123[11], stage122[15], stage121[18], stage120[19]}
   );
   gpc1_1 gpc1_1_2724(
      {stage121[17]},
      {stage121[19]}
   );
   gpc1_1 gpc1_1_2725(
      {stage123[8]},
      {stage123[12]}
   );
   gpc1_1 gpc1_1_2726(
      {stage123[9]},
      {stage123[13]}
   );
   gpc1_1 gpc1_1_2727(
      {stage123[10]},
      {stage123[14]}
   );
   gpc1_1 gpc1_1_2728(
      {stage124[9]},
      {stage124[13]}
   );
   gpc1_1 gpc1_1_2729(
      {stage124[10]},
      {stage124[14]}
   );
   gpc1_1 gpc1_1_2730(
      {stage124[11]},
      {stage124[15]}
   );
   gpc1_1 gpc1_1_2731(
      {stage125[8]},
      {stage125[9]}
   );
   gpc1_1 gpc1_1_2732(
      {stage126[3]},
      {stage126[5]}
   );
   gpc1_1 gpc1_1_2733(
      {stage126[4]},
      {stage126[6]}
   );
   gpc1_1 gpc1_1_2734(
      {stage127[0]},
      {stage127[1]}
   );
   gpc1_1 gpc1_1_2735(
      {stage128[0]},
      {stage128[1]}
   );
   gpc1_1 gpc1_1_2736(
      {stage000[4]},
      {stage000[5]}
   );
   gpc1_1 gpc1_1_2737(
      {stage001[5]},
      {stage001[6]}
   );
   gpc1_1 gpc1_1_2738(
      {stage002[6]},
      {stage002[7]}
   );
   gpc1_1 gpc1_1_2739(
      {stage003[10]},
      {stage003[11]}
   );
   gpc1_1 gpc1_1_2740(
      {stage004[12]},
      {stage004[13]}
   );
   gpc1_1 gpc1_1_2741(
      {stage005[27]},
      {stage005[29]}
   );
   gpc1_1 gpc1_1_2742(
      {stage005[28]},
      {stage005[30]}
   );
   gpc1_1 gpc1_1_2743(
      {stage006[17]},
      {stage006[19]}
   );
   gpc1_1 gpc1_1_2744(
      {stage006[18]},
      {stage006[20]}
   );
   gpc615_5 gpc615_5_2745(
      {stage007[29], stage007[30], stage007[31], stage007[32], stage007[33]},
      {stage008[22]},
      {stage009[36], stage009[37], stage009[38], stage009[39], stage009[40], stage009[41]},
      {stage011[37], stage010[20], stage009[43], stage008[23], stage007[34]}
   );
   gpc1_1 gpc1_1_2746(
      {stage009[42]},
      {stage009[44]}
   );
   gpc1_1 gpc1_1_2747(
      {stage010[19]},
      {stage010[21]}
   );
   gpc135_4 gpc135_4_2748(
      {stage011[32], stage011[33], stage011[34], stage011[35], stage011[36]},
      {stage012[24], stage012[25], 1'h0},
      {stage013[33]},
      {stage014[35], stage013[37], stage012[26], stage011[38]}
   );
   gpc1325_5 gpc1325_5_2749(
      {stage013[34], stage013[35], stage013[36], 1'h0, 1'h0},
      {stage014[34], 1'h0},
      {stage015[36], stage015[37], stage015[38]},
      {stage016[38]},
      {stage017[63], stage016[40], stage015[40], stage014[36], stage013[38]}
   );
   gpc1_1 gpc1_1_2750(
      {stage015[39]},
      {stage015[41]}
   );
   gpc1_1 gpc1_1_2751(
      {stage016[39]},
      {stage016[41]}
   );
   gpc207_4 gpc207_4_2752(
      {stage017[57], stage017[58], stage017[59], stage017[60], stage017[61], stage017[62], 1'h0},
      {stage019[53], 1'h0},
      {stage020[54], stage019[54], stage018[37], stage017[64]}
   );
   gpc1415_5 gpc1415_5_2753(
      {stage018[32], stage018[33], stage018[34], stage018[35], stage018[36]},
      {1'h0},
      {stage020[50], stage020[51], stage020[52], stage020[53]},
      {stage021[48]},
      {stage022[65], stage021[49], stage020[55], stage019[55], stage018[38]}
   );
   gpc615_5 gpc615_5_2754(
      {stage022[60], stage022[61], stage022[62], stage022[63], stage022[64]},
      {stage023[61]},
      {stage024[42], stage024[43], stage024[44], stage024[45], stage024[46], stage024[47]},
      {stage026[64], stage025[68], stage024[48], stage023[63], stage022[66]}
   );
   gpc1_1 gpc1_1_2755(
      {stage023[62]},
      {stage023[64]}
   );
   gpc1_1 gpc1_1_2756(
      {stage025[67]},
      {stage025[69]}
   );
   gpc2135_5 gpc2135_5_2757(
      {stage026[62], stage026[63], 1'h0, 1'h0, 1'h0},
      {stage027[89], stage027[90], stage027[91]},
      {stage028[55]},
      {stage029[66], stage029[67]},
      {stage030[64], stage029[68], stage028[57], stage027[96], stage026[65]}
   );
   gpc15_3 gpc15_3_2758(
      {stage027[92], stage027[93], stage027[94], stage027[95], 1'h0},
      {stage028[56]},
      {stage029[69], stage028[58], stage027[97]}
   );
   gpc207_4 gpc207_4_2759(
      {stage030[61], stage030[62], stage030[63], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage032[94], stage032[95]},
      {stage033[57], stage032[96], stage031[72], stage030[65]}
   );
   gpc207_4 gpc207_4_2760(
      {stage031[65], stage031[66], stage031[67], stage031[68], stage031[69], stage031[70], stage031[71]},
      {stage033[55], stage033[56]},
      {stage034[75], stage033[58], stage032[97], stage031[73]}
   );
   gpc3_2 gpc3_2_2761(
      {stage034[72], stage034[73], stage034[74]},
      {stage035[71], stage034[76]}
   );
   gpc2135_5 gpc2135_5_2762(
      {stage035[66], stage035[67], stage035[68], stage035[69], stage035[70]},
      {stage036[68], stage036[69], stage036[70]},
      {stage037[71]},
      {stage038[89], stage038[90]},
      {stage039[72], stage038[91], stage037[77], stage036[71], stage035[72]}
   );
   gpc606_5 gpc606_5_2763(
      {stage037[72], stage037[73], stage037[74], stage037[75], stage037[76], 1'h0},
      {stage039[66], stage039[67], stage039[68], stage039[69], stage039[70], stage039[71]},
      {stage041[86], stage040[89], stage039[73], stage038[92], stage037[78]}
   );
   gpc2135_5 gpc2135_5_2764(
      {stage040[86], stage040[87], stage040[88], 1'h0, 1'h0},
      {stage041[83], stage041[84], stage041[85]},
      {stage042[89]},
      {stage043[89], stage043[90]},
      {stage044[89], stage043[91], stage042[96], stage041[87], stage040[90]}
   );
   gpc606_5 gpc606_5_2765(
      {stage042[90], stage042[91], stage042[92], stage042[93], stage042[94], stage042[95]},
      {stage044[85], stage044[86], stage044[87], stage044[88], 1'h0, 1'h0},
      {stage046[88], stage045[89], stage044[90], stage043[92], stage042[97]}
   );
   gpc2135_5 gpc2135_5_2766(
      {stage045[84], stage045[85], stage045[86], stage045[87], stage045[88]},
      {stage046[86], stage046[87], 1'h0},
      {stage047[108]},
      {stage048[130], stage048[131]},
      {stage049[100], stage048[133], stage047[112], stage046[89], stage045[90]}
   );
   gpc623_5 gpc623_5_2767(
      {stage047[109], stage047[110], stage047[111]},
      {stage048[132], 1'h0},
      {stage049[94], stage049[95], stage049[96], stage049[97], stage049[98], stage049[99]},
      {stage051[86], stage050[99], stage049[101], stage048[134], stage047[113]}
   );
   gpc223_4 gpc223_4_2768(
      {stage050[96], stage050[97], stage050[98]},
      {stage051[84], stage051[85]},
      {stage052[104], stage052[105]},
      {stage053[138], stage052[107], stage051[87], stage050[100]}
   );
   gpc1_1 gpc1_1_2769(
      {stage052[106]},
      {stage052[108]}
   );
   gpc207_4 gpc207_4_2770(
      {stage053[132], stage053[133], stage053[134], stage053[135], stage053[136], stage053[137], 1'h0},
      {stage055[118], stage055[119]},
      {stage056[101], stage055[122], stage054[128], stage053[139]}
   );
   gpc623_5 gpc623_5_2771(
      {stage054[125], stage054[126], stage054[127]},
      {stage055[120], stage055[121]},
      {stage056[95], stage056[96], stage056[97], stage056[98], stage056[99], stage056[100]},
      {stage058[101], stage057[98], stage056[102], stage055[123], stage054[129]}
   );
   gpc1343_5 gpc1343_5_2772(
      {stage057[95], stage057[96], stage057[97]},
      {stage058[98], stage058[99], stage058[100], 1'h0},
      {stage059[112], stage059[113], stage059[114]},
      {stage060[105]},
      {stage061[135], stage060[107], stage059[116], stage058[102], stage057[99]}
   );
   gpc1_1 gpc1_1_2773(
      {stage059[115]},
      {stage059[117]}
   );
   gpc1_1 gpc1_1_2774(
      {stage060[106]},
      {stage060[108]}
   );
   gpc615_5 gpc615_5_2775(
      {stage061[130], stage061[131], stage061[132], stage061[133], stage061[134]},
      {stage062[135]},
      {stage063[138], stage063[139], stage063[140], stage063[141], stage063[142], stage063[143]},
      {stage065[128], stage064[120], stage063[144], stage062[139], stage061[136]}
   );
   gpc3_2 gpc3_2_2776(
      {stage062[136], stage062[137], stage062[138]},
      {stage063[145], stage062[140]}
   );
   gpc1343_5 gpc1343_5_2777(
      {stage064[117], stage064[118], stage064[119]},
      {stage065[124], stage065[125], stage065[126], stage065[127]},
      {stage066[106], stage066[107], stage066[108]},
      {stage067[121]},
      {stage068[113], stage067[123], stage066[110], stage065[129], stage064[121]}
   );
   gpc1_1 gpc1_1_2778(
      {stage066[109]},
      {stage066[111]}
   );
   gpc1_1 gpc1_1_2779(
      {stage067[122]},
      {stage067[124]}
   );
   gpc207_4 gpc207_4_2780(
      {stage068[107], stage068[108], stage068[109], stage068[110], stage068[111], stage068[112], 1'h0},
      {stage070[108], stage070[109]},
      {stage071[118], stage070[111], stage069[122], stage068[114]}
   );
   gpc615_5 gpc615_5_2781(
      {stage069[117], stage069[118], stage069[119], stage069[120], stage069[121]},
      {stage070[110]},
      {stage071[112], stage071[113], stage071[114], stage071[115], stage071[116], stage071[117]},
      {stage073[101], stage072[110], stage071[119], stage070[112], stage069[123]}
   );
   gpc135_4 gpc135_4_2782(
      {stage072[106], stage072[107], stage072[108], stage072[109], 1'h0},
      {stage073[98], stage073[99], stage073[100]},
      {stage074[114]},
      {stage075[99], stage074[120], stage073[102], stage072[111]}
   );
   gpc2135_5 gpc2135_5_2783(
      {stage074[115], stage074[116], stage074[117], stage074[118], stage074[119]},
      {stage075[96], stage075[97], stage075[98]},
      {stage076[91]},
      {stage077[98], stage077[99]},
      {stage078[101], stage077[102], stage076[95], stage075[100], stage074[121]}
   );
   gpc623_5 gpc623_5_2784(
      {stage076[92], stage076[93], stage076[94]},
      {stage077[100], stage077[101]},
      {stage078[95], stage078[96], stage078[97], stage078[98], stage078[99], stage078[100]},
      {stage080[96], stage079[119], stage078[102], stage077[103], stage076[96]}
   );
   gpc135_4 gpc135_4_2785(
      {stage079[114], stage079[115], stage079[116], stage079[117], stage079[118]},
      {stage080[93], stage080[94], stage080[95]},
      {stage081[95]},
      {stage082[83], stage081[101], stage080[97], stage079[120]}
   );
   gpc2135_5 gpc2135_5_2786(
      {stage081[96], stage081[97], stage081[98], stage081[99], stage081[100]},
      {stage082[80], stage082[81], stage082[82]},
      {stage083[81]},
      {stage084[91], stage084[92]},
      {stage085[88], stage084[93], stage083[88], stage082[84], stage081[102]}
   );
   gpc207_4 gpc207_4_2787(
      {stage083[82], stage083[83], stage083[84], stage083[85], stage083[86], stage083[87], 1'h0},
      {stage085[86], stage085[87]},
      {stage086[87], stage085[89], stage084[94], stage083[89]}
   );
   gpc3_2 gpc3_2_2788(
      {stage086[85], stage086[86], 1'h0},
      {stage087[75], stage086[88]}
   );
   gpc2135_5 gpc2135_5_2789(
      {stage087[71], stage087[72], stage087[73], stage087[74], 1'h0},
      {stage088[73], stage088[74], stage088[75]},
      {stage089[78]},
      {stage090[74], stage090[75]},
      {stage091[87], stage090[78], stage089[82], stage088[77], stage087[76]}
   );
   gpc1_1 gpc1_1_2790(
      {stage088[76]},
      {stage088[78]}
   );
   gpc223_4 gpc223_4_2791(
      {stage089[79], stage089[80], stage089[81]},
      {stage090[76], stage090[77]},
      {stage091[85], stage091[86]},
      {stage092[98], stage091[88], stage090[79], stage089[83]}
   );
   gpc7_3 gpc7_3_2792(
      {stage092[92], stage092[93], stage092[94], stage092[95], stage092[96], stage092[97], 1'h0},
      {stage094[81], stage093[92], stage092[99]}
   );
   gpc2135_5 gpc2135_5_2793(
      {stage093[89], stage093[90], stage093[91], 1'h0, 1'h0},
      {stage094[79], stage094[80], 1'h0},
      {stage095[83]},
      {stage096[57], stage096[58]},
      {stage097[68], stage096[60], stage095[87], stage094[82], stage093[93]}
   );
   gpc615_5 gpc615_5_2794(
      {stage095[84], stage095[85], stage095[86], 1'h0, 1'h0},
      {stage096[59]},
      {stage097[64], stage097[65], stage097[66], stage097[67], 1'h0, 1'h0},
      {stage099[54], stage098[75], stage097[69], stage096[61], stage095[88]}
   );
   gpc2135_5 gpc2135_5_2795(
      {stage098[71], stage098[72], stage098[73], stage098[74], 1'h0},
      {stage099[51], stage099[52], stage099[53]},
      {stage100[61]},
      {stage101[46], stage101[47]},
      {stage102[72], stage101[50], stage100[64], stage099[55], stage098[76]}
   );
   gpc623_5 gpc623_5_2796(
      {stage100[62], stage100[63], 1'h0},
      {stage101[48], stage101[49]},
      {stage102[66], stage102[67], stage102[68], stage102[69], stage102[70], stage102[71]},
      {stage104[39], stage103[58], stage102[73], stage101[51], stage100[65]}
   );
   gpc135_4 gpc135_4_2797(
      {stage103[53], stage103[54], stage103[55], stage103[56], stage103[57]},
      {stage104[38], 1'h0, 1'h0},
      {stage105[76]},
      {stage106[59], stage105[80], stage104[40], stage103[59]}
   );
   gpc1343_5 gpc1343_5_2798(
      {stage105[77], stage105[78], stage105[79]},
      {stage106[55], stage106[56], stage106[57], stage106[58]},
      {stage107[34], stage107[35], 1'h0},
      {stage108[51]},
      {stage109[37], stage108[53], stage107[36], stage106[60], stage105[81]}
   );
   gpc615_5 gpc615_5_2799(
      {1'h0, 1'h0, 1'h0, 1'h0, 1'h0},
      {stage108[52]},
      {stage109[31], stage109[32], stage109[33], stage109[34], stage109[35], stage109[36]},
      {stage111[47], stage110[35], stage109[38], stage108[54], stage107[37]}
   );
   gpc15_3 gpc15_3_2800(
      {stage110[32], stage110[33], stage110[34], 1'h0, 1'h0},
      {stage111[46]},
      {stage112[33], stage111[48], stage110[36]}
   );
   gpc1_1 gpc1_1_2801(
      {stage112[32]},
      {stage112[34]}
   );
   gpc1_1 gpc1_1_2802(
      {stage113[42]},
      {stage113[44]}
   );
   gpc1_1 gpc1_1_2803(
      {stage113[43]},
      {stage113[45]}
   );
   gpc1_1 gpc1_1_2804(
      {stage114[29]},
      {stage114[31]}
   );
   gpc1_1 gpc1_1_2805(
      {stage114[30]},
      {stage114[32]}
   );
   gpc7_3 gpc7_3_2806(
      {stage115[44], stage115[45], stage115[46], stage115[47], 1'h0, 1'h0, 1'h0},
      {stage117[29], stage116[41], stage115[48]}
   );
   gpc23_3 gpc23_3_2807(
      {stage116[39], stage116[40], 1'h0},
      {stage117[27], stage117[28]},
      {stage118[20], stage117[30], stage116[42]}
   );
   gpc15_3 gpc15_3_2808(
      {stage118[17], stage118[18], stage118[19], 1'h0, 1'h0},
      {stage119[25]},
      {stage120[20], stage119[28], stage118[21]}
   );
   gpc15_3 gpc15_3_2809(
      {stage119[26], stage119[27], 1'h0, 1'h0, 1'h0},
      {stage120[19]},
      {stage121[20], stage120[21], stage119[29]}
   );
   gpc615_5 gpc615_5_2810(
      {stage121[18], stage121[19], 1'h0, 1'h0, 1'h0},
      {stage122[15]},
      {stage123[11], stage123[12], stage123[13], stage123[14], 1'h0, 1'h0},
      {stage125[10], stage124[16], stage123[15], stage122[16], stage121[21]}
   );
   gpc215_4 gpc215_4_2811(
      {stage124[12], stage124[13], stage124[14], stage124[15], 1'h0},
      {stage125[9]},
      {stage126[5], stage126[6]},
      {stage127[2], stage126[7], stage125[11], stage124[17]}
   );
   gpc1_1 gpc1_1_2812(
      {stage127[1]},
      {stage127[3]}
   );
   gpc1_1 gpc1_1_2813(
      {stage128[1]},
      {stage128[2]}
   );
endmodule

module behavioral_tester();
   reg [0:0] src000;
   reg [1:0] src001;
   reg [2:0] src002;
   reg [3:0] src003;
   reg [4:0] src004;
   reg [5:0] src005;
   reg [6:0] src006;
   reg [7:0] src007;
   reg [8:0] src008;
   reg [9:0] src009;
   reg [10:0] src010;
   reg [11:0] src011;
   reg [12:0] src012;
   reg [13:0] src013;
   reg [14:0] src014;
   reg [15:0] src015;
   reg [16:0] src016;
   reg [17:0] src017;
   reg [18:0] src018;
   reg [19:0] src019;
   reg [20:0] src020;
   reg [21:0] src021;
   reg [22:0] src022;
   reg [23:0] src023;
   reg [24:0] src024;
   reg [25:0] src025;
   reg [26:0] src026;
   reg [27:0] src027;
   reg [28:0] src028;
   reg [29:0] src029;
   reg [30:0] src030;
   reg [31:0] src031;
   reg [32:0] src032;
   reg [33:0] src033;
   reg [34:0] src034;
   reg [35:0] src035;
   reg [36:0] src036;
   reg [37:0] src037;
   reg [38:0] src038;
   reg [39:0] src039;
   reg [40:0] src040;
   reg [41:0] src041;
   reg [42:0] src042;
   reg [43:0] src043;
   reg [44:0] src044;
   reg [45:0] src045;
   reg [46:0] src046;
   reg [47:0] src047;
   reg [48:0] src048;
   reg [49:0] src049;
   reg [50:0] src050;
   reg [51:0] src051;
   reg [52:0] src052;
   reg [53:0] src053;
   reg [54:0] src054;
   reg [55:0] src055;
   reg [56:0] src056;
   reg [57:0] src057;
   reg [58:0] src058;
   reg [59:0] src059;
   reg [60:0] src060;
   reg [61:0] src061;
   reg [62:0] src062;
   reg [63:0] src063;
   reg [62:0] src064;
   reg [61:0] src065;
   reg [60:0] src066;
   reg [59:0] src067;
   reg [58:0] src068;
   reg [57:0] src069;
   reg [56:0] src070;
   reg [55:0] src071;
   reg [54:0] src072;
   reg [53:0] src073;
   reg [52:0] src074;
   reg [51:0] src075;
   reg [50:0] src076;
   reg [49:0] src077;
   reg [48:0] src078;
   reg [47:0] src079;
   reg [46:0] src080;
   reg [45:0] src081;
   reg [44:0] src082;
   reg [43:0] src083;
   reg [42:0] src084;
   reg [41:0] src085;
   reg [40:0] src086;
   reg [39:0] src087;
   reg [38:0] src088;
   reg [37:0] src089;
   reg [36:0] src090;
   reg [35:0] src091;
   reg [34:0] src092;
   reg [33:0] src093;
   reg [32:0] src094;
   reg [31:0] src095;
   reg [30:0] src096;
   reg [29:0] src097;
   reg [28:0] src098;
   reg [27:0] src099;
   reg [26:0] src100;
   reg [25:0] src101;
   reg [24:0] src102;
   reg [23:0] src103;
   reg [22:0] src104;
   reg [21:0] src105;
   reg [20:0] src106;
   reg [19:0] src107;
   reg [18:0] src108;
   reg [17:0] src109;
   reg [16:0] src110;
   reg [15:0] src111;
   reg [14:0] src112;
   reg [13:0] src113;
   reg [12:0] src114;
   reg [11:0] src115;
   reg [10:0] src116;
   reg [9:0] src117;
   reg [8:0] src118;
   reg [7:0] src119;
   reg [6:0] src120;
   reg [5:0] src121;
   reg [4:0] src122;
   reg [3:0] src123;
   reg [2:0] src124;
   reg [1:0] src125;
   reg [0:0] src126;
   wire [0:0] dst000;
   wire [0:0] dst001;
   wire [0:0] dst002;
   wire [0:0] dst003;
   wire [0:0] dst004;
   wire [1:0] dst005;
   wire [1:0] dst006;
   wire [0:0] dst007;
   wire [0:0] dst008;
   wire [1:0] dst009;
   wire [1:0] dst010;
   wire [1:0] dst011;
   wire [0:0] dst012;
   wire [1:0] dst013;
   wire [1:0] dst014;
   wire [1:0] dst015;
   wire [1:0] dst016;
   wire [1:0] dst017;
   wire [1:0] dst018;
   wire [1:0] dst019;
   wire [1:0] dst020;
   wire [0:0] dst021;
   wire [1:0] dst022;
   wire [1:0] dst023;
   wire [0:0] dst024;
   wire [1:0] dst025;
   wire [1:0] dst026;
   wire [1:0] dst027;
   wire [1:0] dst028;
   wire [1:0] dst029;
   wire [1:0] dst030;
   wire [1:0] dst031;
   wire [1:0] dst032;
   wire [1:0] dst033;
   wire [1:0] dst034;
   wire [1:0] dst035;
   wire [0:0] dst036;
   wire [1:0] dst037;
   wire [1:0] dst038;
   wire [1:0] dst039;
   wire [1:0] dst040;
   wire [1:0] dst041;
   wire [1:0] dst042;
   wire [1:0] dst043;
   wire [1:0] dst044;
   wire [1:0] dst045;
   wire [1:0] dst046;
   wire [1:0] dst047;
   wire [1:0] dst048;
   wire [1:0] dst049;
   wire [1:0] dst050;
   wire [1:0] dst051;
   wire [1:0] dst052;
   wire [1:0] dst053;
   wire [1:0] dst054;
   wire [1:0] dst055;
   wire [1:0] dst056;
   wire [1:0] dst057;
   wire [1:0] dst058;
   wire [1:0] dst059;
   wire [1:0] dst060;
   wire [1:0] dst061;
   wire [1:0] dst062;
   wire [1:0] dst063;
   wire [1:0] dst064;
   wire [1:0] dst065;
   wire [1:0] dst066;
   wire [1:0] dst067;
   wire [1:0] dst068;
   wire [1:0] dst069;
   wire [1:0] dst070;
   wire [1:0] dst071;
   wire [1:0] dst072;
   wire [1:0] dst073;
   wire [1:0] dst074;
   wire [1:0] dst075;
   wire [1:0] dst076;
   wire [1:0] dst077;
   wire [1:0] dst078;
   wire [1:0] dst079;
   wire [1:0] dst080;
   wire [1:0] dst081;
   wire [1:0] dst082;
   wire [1:0] dst083;
   wire [1:0] dst084;
   wire [1:0] dst085;
   wire [1:0] dst086;
   wire [1:0] dst087;
   wire [1:0] dst088;
   wire [1:0] dst089;
   wire [1:0] dst090;
   wire [1:0] dst091;
   wire [1:0] dst092;
   wire [1:0] dst093;
   wire [1:0] dst094;
   wire [1:0] dst095;
   wire [1:0] dst096;
   wire [1:0] dst097;
   wire [1:0] dst098;
   wire [1:0] dst099;
   wire [1:0] dst100;
   wire [1:0] dst101;
   wire [1:0] dst102;
   wire [1:0] dst103;
   wire [1:0] dst104;
   wire [1:0] dst105;
   wire [1:0] dst106;
   wire [1:0] dst107;
   wire [1:0] dst108;
   wire [1:0] dst109;
   wire [1:0] dst110;
   wire [1:0] dst111;
   wire [1:0] dst112;
   wire [1:0] dst113;
   wire [1:0] dst114;
   wire [0:0] dst115;
   wire [1:0] dst116;
   wire [1:0] dst117;
   wire [1:0] dst118;
   wire [1:0] dst119;
   wire [1:0] dst120;
   wire [1:0] dst121;
   wire [0:0] dst122;
   wire [0:0] dst123;
   wire [1:0] dst124;
   wire [1:0] dst125;
   wire [0:0] dst126;
   wire [1:0] dst127;
   wire [0:0] dst128;
   wire [129:0] srcsum;
   wire [129:0] dstsum;
   wire test;
   assign srcsum =
      (src000[0] << 0) +
      (src001[0] << 1) +
      (src001[1] << 1) +
      (src002[0] << 2) +
      (src002[1] << 2) +
      (src002[2] << 2) +
      (src003[0] << 3) +
      (src003[1] << 3) +
      (src003[2] << 3) +
      (src003[3] << 3) +
      (src004[0] << 4) +
      (src004[1] << 4) +
      (src004[2] << 4) +
      (src004[3] << 4) +
      (src004[4] << 4) +
      (src005[0] << 5) +
      (src005[1] << 5) +
      (src005[2] << 5) +
      (src005[3] << 5) +
      (src005[4] << 5) +
      (src005[5] << 5) +
      (src006[0] << 6) +
      (src006[1] << 6) +
      (src006[2] << 6) +
      (src006[3] << 6) +
      (src006[4] << 6) +
      (src006[5] << 6) +
      (src006[6] << 6) +
      (src007[0] << 7) +
      (src007[1] << 7) +
      (src007[2] << 7) +
      (src007[3] << 7) +
      (src007[4] << 7) +
      (src007[5] << 7) +
      (src007[6] << 7) +
      (src007[7] << 7) +
      (src008[0] << 8) +
      (src008[1] << 8) +
      (src008[2] << 8) +
      (src008[3] << 8) +
      (src008[4] << 8) +
      (src008[5] << 8) +
      (src008[6] << 8) +
      (src008[7] << 8) +
      (src008[8] << 8) +
      (src009[0] << 9) +
      (src009[1] << 9) +
      (src009[2] << 9) +
      (src009[3] << 9) +
      (src009[4] << 9) +
      (src009[5] << 9) +
      (src009[6] << 9) +
      (src009[7] << 9) +
      (src009[8] << 9) +
      (src009[9] << 9) +
      (src010[0] << 10) +
      (src010[1] << 10) +
      (src010[2] << 10) +
      (src010[3] << 10) +
      (src010[4] << 10) +
      (src010[5] << 10) +
      (src010[6] << 10) +
      (src010[7] << 10) +
      (src010[8] << 10) +
      (src010[9] << 10) +
      (src010[10] << 10) +
      (src011[0] << 11) +
      (src011[1] << 11) +
      (src011[2] << 11) +
      (src011[3] << 11) +
      (src011[4] << 11) +
      (src011[5] << 11) +
      (src011[6] << 11) +
      (src011[7] << 11) +
      (src011[8] << 11) +
      (src011[9] << 11) +
      (src011[10] << 11) +
      (src011[11] << 11) +
      (src012[0] << 12) +
      (src012[1] << 12) +
      (src012[2] << 12) +
      (src012[3] << 12) +
      (src012[4] << 12) +
      (src012[5] << 12) +
      (src012[6] << 12) +
      (src012[7] << 12) +
      (src012[8] << 12) +
      (src012[9] << 12) +
      (src012[10] << 12) +
      (src012[11] << 12) +
      (src012[12] << 12) +
      (src013[0] << 13) +
      (src013[1] << 13) +
      (src013[2] << 13) +
      (src013[3] << 13) +
      (src013[4] << 13) +
      (src013[5] << 13) +
      (src013[6] << 13) +
      (src013[7] << 13) +
      (src013[8] << 13) +
      (src013[9] << 13) +
      (src013[10] << 13) +
      (src013[11] << 13) +
      (src013[12] << 13) +
      (src013[13] << 13) +
      (src014[0] << 14) +
      (src014[1] << 14) +
      (src014[2] << 14) +
      (src014[3] << 14) +
      (src014[4] << 14) +
      (src014[5] << 14) +
      (src014[6] << 14) +
      (src014[7] << 14) +
      (src014[8] << 14) +
      (src014[9] << 14) +
      (src014[10] << 14) +
      (src014[11] << 14) +
      (src014[12] << 14) +
      (src014[13] << 14) +
      (src014[14] << 14) +
      (src015[0] << 15) +
      (src015[1] << 15) +
      (src015[2] << 15) +
      (src015[3] << 15) +
      (src015[4] << 15) +
      (src015[5] << 15) +
      (src015[6] << 15) +
      (src015[7] << 15) +
      (src015[8] << 15) +
      (src015[9] << 15) +
      (src015[10] << 15) +
      (src015[11] << 15) +
      (src015[12] << 15) +
      (src015[13] << 15) +
      (src015[14] << 15) +
      (src015[15] << 15) +
      (src016[0] << 16) +
      (src016[1] << 16) +
      (src016[2] << 16) +
      (src016[3] << 16) +
      (src016[4] << 16) +
      (src016[5] << 16) +
      (src016[6] << 16) +
      (src016[7] << 16) +
      (src016[8] << 16) +
      (src016[9] << 16) +
      (src016[10] << 16) +
      (src016[11] << 16) +
      (src016[12] << 16) +
      (src016[13] << 16) +
      (src016[14] << 16) +
      (src016[15] << 16) +
      (src016[16] << 16) +
      (src017[0] << 17) +
      (src017[1] << 17) +
      (src017[2] << 17) +
      (src017[3] << 17) +
      (src017[4] << 17) +
      (src017[5] << 17) +
      (src017[6] << 17) +
      (src017[7] << 17) +
      (src017[8] << 17) +
      (src017[9] << 17) +
      (src017[10] << 17) +
      (src017[11] << 17) +
      (src017[12] << 17) +
      (src017[13] << 17) +
      (src017[14] << 17) +
      (src017[15] << 17) +
      (src017[16] << 17) +
      (src017[17] << 17) +
      (src018[0] << 18) +
      (src018[1] << 18) +
      (src018[2] << 18) +
      (src018[3] << 18) +
      (src018[4] << 18) +
      (src018[5] << 18) +
      (src018[6] << 18) +
      (src018[7] << 18) +
      (src018[8] << 18) +
      (src018[9] << 18) +
      (src018[10] << 18) +
      (src018[11] << 18) +
      (src018[12] << 18) +
      (src018[13] << 18) +
      (src018[14] << 18) +
      (src018[15] << 18) +
      (src018[16] << 18) +
      (src018[17] << 18) +
      (src018[18] << 18) +
      (src019[0] << 19) +
      (src019[1] << 19) +
      (src019[2] << 19) +
      (src019[3] << 19) +
      (src019[4] << 19) +
      (src019[5] << 19) +
      (src019[6] << 19) +
      (src019[7] << 19) +
      (src019[8] << 19) +
      (src019[9] << 19) +
      (src019[10] << 19) +
      (src019[11] << 19) +
      (src019[12] << 19) +
      (src019[13] << 19) +
      (src019[14] << 19) +
      (src019[15] << 19) +
      (src019[16] << 19) +
      (src019[17] << 19) +
      (src019[18] << 19) +
      (src019[19] << 19) +
      (src020[0] << 20) +
      (src020[1] << 20) +
      (src020[2] << 20) +
      (src020[3] << 20) +
      (src020[4] << 20) +
      (src020[5] << 20) +
      (src020[6] << 20) +
      (src020[7] << 20) +
      (src020[8] << 20) +
      (src020[9] << 20) +
      (src020[10] << 20) +
      (src020[11] << 20) +
      (src020[12] << 20) +
      (src020[13] << 20) +
      (src020[14] << 20) +
      (src020[15] << 20) +
      (src020[16] << 20) +
      (src020[17] << 20) +
      (src020[18] << 20) +
      (src020[19] << 20) +
      (src020[20] << 20) +
      (src021[0] << 21) +
      (src021[1] << 21) +
      (src021[2] << 21) +
      (src021[3] << 21) +
      (src021[4] << 21) +
      (src021[5] << 21) +
      (src021[6] << 21) +
      (src021[7] << 21) +
      (src021[8] << 21) +
      (src021[9] << 21) +
      (src021[10] << 21) +
      (src021[11] << 21) +
      (src021[12] << 21) +
      (src021[13] << 21) +
      (src021[14] << 21) +
      (src021[15] << 21) +
      (src021[16] << 21) +
      (src021[17] << 21) +
      (src021[18] << 21) +
      (src021[19] << 21) +
      (src021[20] << 21) +
      (src021[21] << 21) +
      (src022[0] << 22) +
      (src022[1] << 22) +
      (src022[2] << 22) +
      (src022[3] << 22) +
      (src022[4] << 22) +
      (src022[5] << 22) +
      (src022[6] << 22) +
      (src022[7] << 22) +
      (src022[8] << 22) +
      (src022[9] << 22) +
      (src022[10] << 22) +
      (src022[11] << 22) +
      (src022[12] << 22) +
      (src022[13] << 22) +
      (src022[14] << 22) +
      (src022[15] << 22) +
      (src022[16] << 22) +
      (src022[17] << 22) +
      (src022[18] << 22) +
      (src022[19] << 22) +
      (src022[20] << 22) +
      (src022[21] << 22) +
      (src022[22] << 22) +
      (src023[0] << 23) +
      (src023[1] << 23) +
      (src023[2] << 23) +
      (src023[3] << 23) +
      (src023[4] << 23) +
      (src023[5] << 23) +
      (src023[6] << 23) +
      (src023[7] << 23) +
      (src023[8] << 23) +
      (src023[9] << 23) +
      (src023[10] << 23) +
      (src023[11] << 23) +
      (src023[12] << 23) +
      (src023[13] << 23) +
      (src023[14] << 23) +
      (src023[15] << 23) +
      (src023[16] << 23) +
      (src023[17] << 23) +
      (src023[18] << 23) +
      (src023[19] << 23) +
      (src023[20] << 23) +
      (src023[21] << 23) +
      (src023[22] << 23) +
      (src023[23] << 23) +
      (src024[0] << 24) +
      (src024[1] << 24) +
      (src024[2] << 24) +
      (src024[3] << 24) +
      (src024[4] << 24) +
      (src024[5] << 24) +
      (src024[6] << 24) +
      (src024[7] << 24) +
      (src024[8] << 24) +
      (src024[9] << 24) +
      (src024[10] << 24) +
      (src024[11] << 24) +
      (src024[12] << 24) +
      (src024[13] << 24) +
      (src024[14] << 24) +
      (src024[15] << 24) +
      (src024[16] << 24) +
      (src024[17] << 24) +
      (src024[18] << 24) +
      (src024[19] << 24) +
      (src024[20] << 24) +
      (src024[21] << 24) +
      (src024[22] << 24) +
      (src024[23] << 24) +
      (src024[24] << 24) +
      (src025[0] << 25) +
      (src025[1] << 25) +
      (src025[2] << 25) +
      (src025[3] << 25) +
      (src025[4] << 25) +
      (src025[5] << 25) +
      (src025[6] << 25) +
      (src025[7] << 25) +
      (src025[8] << 25) +
      (src025[9] << 25) +
      (src025[10] << 25) +
      (src025[11] << 25) +
      (src025[12] << 25) +
      (src025[13] << 25) +
      (src025[14] << 25) +
      (src025[15] << 25) +
      (src025[16] << 25) +
      (src025[17] << 25) +
      (src025[18] << 25) +
      (src025[19] << 25) +
      (src025[20] << 25) +
      (src025[21] << 25) +
      (src025[22] << 25) +
      (src025[23] << 25) +
      (src025[24] << 25) +
      (src025[25] << 25) +
      (src026[0] << 26) +
      (src026[1] << 26) +
      (src026[2] << 26) +
      (src026[3] << 26) +
      (src026[4] << 26) +
      (src026[5] << 26) +
      (src026[6] << 26) +
      (src026[7] << 26) +
      (src026[8] << 26) +
      (src026[9] << 26) +
      (src026[10] << 26) +
      (src026[11] << 26) +
      (src026[12] << 26) +
      (src026[13] << 26) +
      (src026[14] << 26) +
      (src026[15] << 26) +
      (src026[16] << 26) +
      (src026[17] << 26) +
      (src026[18] << 26) +
      (src026[19] << 26) +
      (src026[20] << 26) +
      (src026[21] << 26) +
      (src026[22] << 26) +
      (src026[23] << 26) +
      (src026[24] << 26) +
      (src026[25] << 26) +
      (src026[26] << 26) +
      (src027[0] << 27) +
      (src027[1] << 27) +
      (src027[2] << 27) +
      (src027[3] << 27) +
      (src027[4] << 27) +
      (src027[5] << 27) +
      (src027[6] << 27) +
      (src027[7] << 27) +
      (src027[8] << 27) +
      (src027[9] << 27) +
      (src027[10] << 27) +
      (src027[11] << 27) +
      (src027[12] << 27) +
      (src027[13] << 27) +
      (src027[14] << 27) +
      (src027[15] << 27) +
      (src027[16] << 27) +
      (src027[17] << 27) +
      (src027[18] << 27) +
      (src027[19] << 27) +
      (src027[20] << 27) +
      (src027[21] << 27) +
      (src027[22] << 27) +
      (src027[23] << 27) +
      (src027[24] << 27) +
      (src027[25] << 27) +
      (src027[26] << 27) +
      (src027[27] << 27) +
      (src028[0] << 28) +
      (src028[1] << 28) +
      (src028[2] << 28) +
      (src028[3] << 28) +
      (src028[4] << 28) +
      (src028[5] << 28) +
      (src028[6] << 28) +
      (src028[7] << 28) +
      (src028[8] << 28) +
      (src028[9] << 28) +
      (src028[10] << 28) +
      (src028[11] << 28) +
      (src028[12] << 28) +
      (src028[13] << 28) +
      (src028[14] << 28) +
      (src028[15] << 28) +
      (src028[16] << 28) +
      (src028[17] << 28) +
      (src028[18] << 28) +
      (src028[19] << 28) +
      (src028[20] << 28) +
      (src028[21] << 28) +
      (src028[22] << 28) +
      (src028[23] << 28) +
      (src028[24] << 28) +
      (src028[25] << 28) +
      (src028[26] << 28) +
      (src028[27] << 28) +
      (src028[28] << 28) +
      (src029[0] << 29) +
      (src029[1] << 29) +
      (src029[2] << 29) +
      (src029[3] << 29) +
      (src029[4] << 29) +
      (src029[5] << 29) +
      (src029[6] << 29) +
      (src029[7] << 29) +
      (src029[8] << 29) +
      (src029[9] << 29) +
      (src029[10] << 29) +
      (src029[11] << 29) +
      (src029[12] << 29) +
      (src029[13] << 29) +
      (src029[14] << 29) +
      (src029[15] << 29) +
      (src029[16] << 29) +
      (src029[17] << 29) +
      (src029[18] << 29) +
      (src029[19] << 29) +
      (src029[20] << 29) +
      (src029[21] << 29) +
      (src029[22] << 29) +
      (src029[23] << 29) +
      (src029[24] << 29) +
      (src029[25] << 29) +
      (src029[26] << 29) +
      (src029[27] << 29) +
      (src029[28] << 29) +
      (src029[29] << 29) +
      (src030[0] << 30) +
      (src030[1] << 30) +
      (src030[2] << 30) +
      (src030[3] << 30) +
      (src030[4] << 30) +
      (src030[5] << 30) +
      (src030[6] << 30) +
      (src030[7] << 30) +
      (src030[8] << 30) +
      (src030[9] << 30) +
      (src030[10] << 30) +
      (src030[11] << 30) +
      (src030[12] << 30) +
      (src030[13] << 30) +
      (src030[14] << 30) +
      (src030[15] << 30) +
      (src030[16] << 30) +
      (src030[17] << 30) +
      (src030[18] << 30) +
      (src030[19] << 30) +
      (src030[20] << 30) +
      (src030[21] << 30) +
      (src030[22] << 30) +
      (src030[23] << 30) +
      (src030[24] << 30) +
      (src030[25] << 30) +
      (src030[26] << 30) +
      (src030[27] << 30) +
      (src030[28] << 30) +
      (src030[29] << 30) +
      (src030[30] << 30) +
      (src031[0] << 31) +
      (src031[1] << 31) +
      (src031[2] << 31) +
      (src031[3] << 31) +
      (src031[4] << 31) +
      (src031[5] << 31) +
      (src031[6] << 31) +
      (src031[7] << 31) +
      (src031[8] << 31) +
      (src031[9] << 31) +
      (src031[10] << 31) +
      (src031[11] << 31) +
      (src031[12] << 31) +
      (src031[13] << 31) +
      (src031[14] << 31) +
      (src031[15] << 31) +
      (src031[16] << 31) +
      (src031[17] << 31) +
      (src031[18] << 31) +
      (src031[19] << 31) +
      (src031[20] << 31) +
      (src031[21] << 31) +
      (src031[22] << 31) +
      (src031[23] << 31) +
      (src031[24] << 31) +
      (src031[25] << 31) +
      (src031[26] << 31) +
      (src031[27] << 31) +
      (src031[28] << 31) +
      (src031[29] << 31) +
      (src031[30] << 31) +
      (src031[31] << 31) +
      (src032[0] << 32) +
      (src032[1] << 32) +
      (src032[2] << 32) +
      (src032[3] << 32) +
      (src032[4] << 32) +
      (src032[5] << 32) +
      (src032[6] << 32) +
      (src032[7] << 32) +
      (src032[8] << 32) +
      (src032[9] << 32) +
      (src032[10] << 32) +
      (src032[11] << 32) +
      (src032[12] << 32) +
      (src032[13] << 32) +
      (src032[14] << 32) +
      (src032[15] << 32) +
      (src032[16] << 32) +
      (src032[17] << 32) +
      (src032[18] << 32) +
      (src032[19] << 32) +
      (src032[20] << 32) +
      (src032[21] << 32) +
      (src032[22] << 32) +
      (src032[23] << 32) +
      (src032[24] << 32) +
      (src032[25] << 32) +
      (src032[26] << 32) +
      (src032[27] << 32) +
      (src032[28] << 32) +
      (src032[29] << 32) +
      (src032[30] << 32) +
      (src032[31] << 32) +
      (src032[32] << 32) +
      (src033[0] << 33) +
      (src033[1] << 33) +
      (src033[2] << 33) +
      (src033[3] << 33) +
      (src033[4] << 33) +
      (src033[5] << 33) +
      (src033[6] << 33) +
      (src033[7] << 33) +
      (src033[8] << 33) +
      (src033[9] << 33) +
      (src033[10] << 33) +
      (src033[11] << 33) +
      (src033[12] << 33) +
      (src033[13] << 33) +
      (src033[14] << 33) +
      (src033[15] << 33) +
      (src033[16] << 33) +
      (src033[17] << 33) +
      (src033[18] << 33) +
      (src033[19] << 33) +
      (src033[20] << 33) +
      (src033[21] << 33) +
      (src033[22] << 33) +
      (src033[23] << 33) +
      (src033[24] << 33) +
      (src033[25] << 33) +
      (src033[26] << 33) +
      (src033[27] << 33) +
      (src033[28] << 33) +
      (src033[29] << 33) +
      (src033[30] << 33) +
      (src033[31] << 33) +
      (src033[32] << 33) +
      (src033[33] << 33) +
      (src034[0] << 34) +
      (src034[1] << 34) +
      (src034[2] << 34) +
      (src034[3] << 34) +
      (src034[4] << 34) +
      (src034[5] << 34) +
      (src034[6] << 34) +
      (src034[7] << 34) +
      (src034[8] << 34) +
      (src034[9] << 34) +
      (src034[10] << 34) +
      (src034[11] << 34) +
      (src034[12] << 34) +
      (src034[13] << 34) +
      (src034[14] << 34) +
      (src034[15] << 34) +
      (src034[16] << 34) +
      (src034[17] << 34) +
      (src034[18] << 34) +
      (src034[19] << 34) +
      (src034[20] << 34) +
      (src034[21] << 34) +
      (src034[22] << 34) +
      (src034[23] << 34) +
      (src034[24] << 34) +
      (src034[25] << 34) +
      (src034[26] << 34) +
      (src034[27] << 34) +
      (src034[28] << 34) +
      (src034[29] << 34) +
      (src034[30] << 34) +
      (src034[31] << 34) +
      (src034[32] << 34) +
      (src034[33] << 34) +
      (src034[34] << 34) +
      (src035[0] << 35) +
      (src035[1] << 35) +
      (src035[2] << 35) +
      (src035[3] << 35) +
      (src035[4] << 35) +
      (src035[5] << 35) +
      (src035[6] << 35) +
      (src035[7] << 35) +
      (src035[8] << 35) +
      (src035[9] << 35) +
      (src035[10] << 35) +
      (src035[11] << 35) +
      (src035[12] << 35) +
      (src035[13] << 35) +
      (src035[14] << 35) +
      (src035[15] << 35) +
      (src035[16] << 35) +
      (src035[17] << 35) +
      (src035[18] << 35) +
      (src035[19] << 35) +
      (src035[20] << 35) +
      (src035[21] << 35) +
      (src035[22] << 35) +
      (src035[23] << 35) +
      (src035[24] << 35) +
      (src035[25] << 35) +
      (src035[26] << 35) +
      (src035[27] << 35) +
      (src035[28] << 35) +
      (src035[29] << 35) +
      (src035[30] << 35) +
      (src035[31] << 35) +
      (src035[32] << 35) +
      (src035[33] << 35) +
      (src035[34] << 35) +
      (src035[35] << 35) +
      (src036[0] << 36) +
      (src036[1] << 36) +
      (src036[2] << 36) +
      (src036[3] << 36) +
      (src036[4] << 36) +
      (src036[5] << 36) +
      (src036[6] << 36) +
      (src036[7] << 36) +
      (src036[8] << 36) +
      (src036[9] << 36) +
      (src036[10] << 36) +
      (src036[11] << 36) +
      (src036[12] << 36) +
      (src036[13] << 36) +
      (src036[14] << 36) +
      (src036[15] << 36) +
      (src036[16] << 36) +
      (src036[17] << 36) +
      (src036[18] << 36) +
      (src036[19] << 36) +
      (src036[20] << 36) +
      (src036[21] << 36) +
      (src036[22] << 36) +
      (src036[23] << 36) +
      (src036[24] << 36) +
      (src036[25] << 36) +
      (src036[26] << 36) +
      (src036[27] << 36) +
      (src036[28] << 36) +
      (src036[29] << 36) +
      (src036[30] << 36) +
      (src036[31] << 36) +
      (src036[32] << 36) +
      (src036[33] << 36) +
      (src036[34] << 36) +
      (src036[35] << 36) +
      (src036[36] << 36) +
      (src037[0] << 37) +
      (src037[1] << 37) +
      (src037[2] << 37) +
      (src037[3] << 37) +
      (src037[4] << 37) +
      (src037[5] << 37) +
      (src037[6] << 37) +
      (src037[7] << 37) +
      (src037[8] << 37) +
      (src037[9] << 37) +
      (src037[10] << 37) +
      (src037[11] << 37) +
      (src037[12] << 37) +
      (src037[13] << 37) +
      (src037[14] << 37) +
      (src037[15] << 37) +
      (src037[16] << 37) +
      (src037[17] << 37) +
      (src037[18] << 37) +
      (src037[19] << 37) +
      (src037[20] << 37) +
      (src037[21] << 37) +
      (src037[22] << 37) +
      (src037[23] << 37) +
      (src037[24] << 37) +
      (src037[25] << 37) +
      (src037[26] << 37) +
      (src037[27] << 37) +
      (src037[28] << 37) +
      (src037[29] << 37) +
      (src037[30] << 37) +
      (src037[31] << 37) +
      (src037[32] << 37) +
      (src037[33] << 37) +
      (src037[34] << 37) +
      (src037[35] << 37) +
      (src037[36] << 37) +
      (src037[37] << 37) +
      (src038[0] << 38) +
      (src038[1] << 38) +
      (src038[2] << 38) +
      (src038[3] << 38) +
      (src038[4] << 38) +
      (src038[5] << 38) +
      (src038[6] << 38) +
      (src038[7] << 38) +
      (src038[8] << 38) +
      (src038[9] << 38) +
      (src038[10] << 38) +
      (src038[11] << 38) +
      (src038[12] << 38) +
      (src038[13] << 38) +
      (src038[14] << 38) +
      (src038[15] << 38) +
      (src038[16] << 38) +
      (src038[17] << 38) +
      (src038[18] << 38) +
      (src038[19] << 38) +
      (src038[20] << 38) +
      (src038[21] << 38) +
      (src038[22] << 38) +
      (src038[23] << 38) +
      (src038[24] << 38) +
      (src038[25] << 38) +
      (src038[26] << 38) +
      (src038[27] << 38) +
      (src038[28] << 38) +
      (src038[29] << 38) +
      (src038[30] << 38) +
      (src038[31] << 38) +
      (src038[32] << 38) +
      (src038[33] << 38) +
      (src038[34] << 38) +
      (src038[35] << 38) +
      (src038[36] << 38) +
      (src038[37] << 38) +
      (src038[38] << 38) +
      (src039[0] << 39) +
      (src039[1] << 39) +
      (src039[2] << 39) +
      (src039[3] << 39) +
      (src039[4] << 39) +
      (src039[5] << 39) +
      (src039[6] << 39) +
      (src039[7] << 39) +
      (src039[8] << 39) +
      (src039[9] << 39) +
      (src039[10] << 39) +
      (src039[11] << 39) +
      (src039[12] << 39) +
      (src039[13] << 39) +
      (src039[14] << 39) +
      (src039[15] << 39) +
      (src039[16] << 39) +
      (src039[17] << 39) +
      (src039[18] << 39) +
      (src039[19] << 39) +
      (src039[20] << 39) +
      (src039[21] << 39) +
      (src039[22] << 39) +
      (src039[23] << 39) +
      (src039[24] << 39) +
      (src039[25] << 39) +
      (src039[26] << 39) +
      (src039[27] << 39) +
      (src039[28] << 39) +
      (src039[29] << 39) +
      (src039[30] << 39) +
      (src039[31] << 39) +
      (src039[32] << 39) +
      (src039[33] << 39) +
      (src039[34] << 39) +
      (src039[35] << 39) +
      (src039[36] << 39) +
      (src039[37] << 39) +
      (src039[38] << 39) +
      (src039[39] << 39) +
      (src040[0] << 40) +
      (src040[1] << 40) +
      (src040[2] << 40) +
      (src040[3] << 40) +
      (src040[4] << 40) +
      (src040[5] << 40) +
      (src040[6] << 40) +
      (src040[7] << 40) +
      (src040[8] << 40) +
      (src040[9] << 40) +
      (src040[10] << 40) +
      (src040[11] << 40) +
      (src040[12] << 40) +
      (src040[13] << 40) +
      (src040[14] << 40) +
      (src040[15] << 40) +
      (src040[16] << 40) +
      (src040[17] << 40) +
      (src040[18] << 40) +
      (src040[19] << 40) +
      (src040[20] << 40) +
      (src040[21] << 40) +
      (src040[22] << 40) +
      (src040[23] << 40) +
      (src040[24] << 40) +
      (src040[25] << 40) +
      (src040[26] << 40) +
      (src040[27] << 40) +
      (src040[28] << 40) +
      (src040[29] << 40) +
      (src040[30] << 40) +
      (src040[31] << 40) +
      (src040[32] << 40) +
      (src040[33] << 40) +
      (src040[34] << 40) +
      (src040[35] << 40) +
      (src040[36] << 40) +
      (src040[37] << 40) +
      (src040[38] << 40) +
      (src040[39] << 40) +
      (src040[40] << 40) +
      (src041[0] << 41) +
      (src041[1] << 41) +
      (src041[2] << 41) +
      (src041[3] << 41) +
      (src041[4] << 41) +
      (src041[5] << 41) +
      (src041[6] << 41) +
      (src041[7] << 41) +
      (src041[8] << 41) +
      (src041[9] << 41) +
      (src041[10] << 41) +
      (src041[11] << 41) +
      (src041[12] << 41) +
      (src041[13] << 41) +
      (src041[14] << 41) +
      (src041[15] << 41) +
      (src041[16] << 41) +
      (src041[17] << 41) +
      (src041[18] << 41) +
      (src041[19] << 41) +
      (src041[20] << 41) +
      (src041[21] << 41) +
      (src041[22] << 41) +
      (src041[23] << 41) +
      (src041[24] << 41) +
      (src041[25] << 41) +
      (src041[26] << 41) +
      (src041[27] << 41) +
      (src041[28] << 41) +
      (src041[29] << 41) +
      (src041[30] << 41) +
      (src041[31] << 41) +
      (src041[32] << 41) +
      (src041[33] << 41) +
      (src041[34] << 41) +
      (src041[35] << 41) +
      (src041[36] << 41) +
      (src041[37] << 41) +
      (src041[38] << 41) +
      (src041[39] << 41) +
      (src041[40] << 41) +
      (src041[41] << 41) +
      (src042[0] << 42) +
      (src042[1] << 42) +
      (src042[2] << 42) +
      (src042[3] << 42) +
      (src042[4] << 42) +
      (src042[5] << 42) +
      (src042[6] << 42) +
      (src042[7] << 42) +
      (src042[8] << 42) +
      (src042[9] << 42) +
      (src042[10] << 42) +
      (src042[11] << 42) +
      (src042[12] << 42) +
      (src042[13] << 42) +
      (src042[14] << 42) +
      (src042[15] << 42) +
      (src042[16] << 42) +
      (src042[17] << 42) +
      (src042[18] << 42) +
      (src042[19] << 42) +
      (src042[20] << 42) +
      (src042[21] << 42) +
      (src042[22] << 42) +
      (src042[23] << 42) +
      (src042[24] << 42) +
      (src042[25] << 42) +
      (src042[26] << 42) +
      (src042[27] << 42) +
      (src042[28] << 42) +
      (src042[29] << 42) +
      (src042[30] << 42) +
      (src042[31] << 42) +
      (src042[32] << 42) +
      (src042[33] << 42) +
      (src042[34] << 42) +
      (src042[35] << 42) +
      (src042[36] << 42) +
      (src042[37] << 42) +
      (src042[38] << 42) +
      (src042[39] << 42) +
      (src042[40] << 42) +
      (src042[41] << 42) +
      (src042[42] << 42) +
      (src043[0] << 43) +
      (src043[1] << 43) +
      (src043[2] << 43) +
      (src043[3] << 43) +
      (src043[4] << 43) +
      (src043[5] << 43) +
      (src043[6] << 43) +
      (src043[7] << 43) +
      (src043[8] << 43) +
      (src043[9] << 43) +
      (src043[10] << 43) +
      (src043[11] << 43) +
      (src043[12] << 43) +
      (src043[13] << 43) +
      (src043[14] << 43) +
      (src043[15] << 43) +
      (src043[16] << 43) +
      (src043[17] << 43) +
      (src043[18] << 43) +
      (src043[19] << 43) +
      (src043[20] << 43) +
      (src043[21] << 43) +
      (src043[22] << 43) +
      (src043[23] << 43) +
      (src043[24] << 43) +
      (src043[25] << 43) +
      (src043[26] << 43) +
      (src043[27] << 43) +
      (src043[28] << 43) +
      (src043[29] << 43) +
      (src043[30] << 43) +
      (src043[31] << 43) +
      (src043[32] << 43) +
      (src043[33] << 43) +
      (src043[34] << 43) +
      (src043[35] << 43) +
      (src043[36] << 43) +
      (src043[37] << 43) +
      (src043[38] << 43) +
      (src043[39] << 43) +
      (src043[40] << 43) +
      (src043[41] << 43) +
      (src043[42] << 43) +
      (src043[43] << 43) +
      (src044[0] << 44) +
      (src044[1] << 44) +
      (src044[2] << 44) +
      (src044[3] << 44) +
      (src044[4] << 44) +
      (src044[5] << 44) +
      (src044[6] << 44) +
      (src044[7] << 44) +
      (src044[8] << 44) +
      (src044[9] << 44) +
      (src044[10] << 44) +
      (src044[11] << 44) +
      (src044[12] << 44) +
      (src044[13] << 44) +
      (src044[14] << 44) +
      (src044[15] << 44) +
      (src044[16] << 44) +
      (src044[17] << 44) +
      (src044[18] << 44) +
      (src044[19] << 44) +
      (src044[20] << 44) +
      (src044[21] << 44) +
      (src044[22] << 44) +
      (src044[23] << 44) +
      (src044[24] << 44) +
      (src044[25] << 44) +
      (src044[26] << 44) +
      (src044[27] << 44) +
      (src044[28] << 44) +
      (src044[29] << 44) +
      (src044[30] << 44) +
      (src044[31] << 44) +
      (src044[32] << 44) +
      (src044[33] << 44) +
      (src044[34] << 44) +
      (src044[35] << 44) +
      (src044[36] << 44) +
      (src044[37] << 44) +
      (src044[38] << 44) +
      (src044[39] << 44) +
      (src044[40] << 44) +
      (src044[41] << 44) +
      (src044[42] << 44) +
      (src044[43] << 44) +
      (src044[44] << 44) +
      (src045[0] << 45) +
      (src045[1] << 45) +
      (src045[2] << 45) +
      (src045[3] << 45) +
      (src045[4] << 45) +
      (src045[5] << 45) +
      (src045[6] << 45) +
      (src045[7] << 45) +
      (src045[8] << 45) +
      (src045[9] << 45) +
      (src045[10] << 45) +
      (src045[11] << 45) +
      (src045[12] << 45) +
      (src045[13] << 45) +
      (src045[14] << 45) +
      (src045[15] << 45) +
      (src045[16] << 45) +
      (src045[17] << 45) +
      (src045[18] << 45) +
      (src045[19] << 45) +
      (src045[20] << 45) +
      (src045[21] << 45) +
      (src045[22] << 45) +
      (src045[23] << 45) +
      (src045[24] << 45) +
      (src045[25] << 45) +
      (src045[26] << 45) +
      (src045[27] << 45) +
      (src045[28] << 45) +
      (src045[29] << 45) +
      (src045[30] << 45) +
      (src045[31] << 45) +
      (src045[32] << 45) +
      (src045[33] << 45) +
      (src045[34] << 45) +
      (src045[35] << 45) +
      (src045[36] << 45) +
      (src045[37] << 45) +
      (src045[38] << 45) +
      (src045[39] << 45) +
      (src045[40] << 45) +
      (src045[41] << 45) +
      (src045[42] << 45) +
      (src045[43] << 45) +
      (src045[44] << 45) +
      (src045[45] << 45) +
      (src046[0] << 46) +
      (src046[1] << 46) +
      (src046[2] << 46) +
      (src046[3] << 46) +
      (src046[4] << 46) +
      (src046[5] << 46) +
      (src046[6] << 46) +
      (src046[7] << 46) +
      (src046[8] << 46) +
      (src046[9] << 46) +
      (src046[10] << 46) +
      (src046[11] << 46) +
      (src046[12] << 46) +
      (src046[13] << 46) +
      (src046[14] << 46) +
      (src046[15] << 46) +
      (src046[16] << 46) +
      (src046[17] << 46) +
      (src046[18] << 46) +
      (src046[19] << 46) +
      (src046[20] << 46) +
      (src046[21] << 46) +
      (src046[22] << 46) +
      (src046[23] << 46) +
      (src046[24] << 46) +
      (src046[25] << 46) +
      (src046[26] << 46) +
      (src046[27] << 46) +
      (src046[28] << 46) +
      (src046[29] << 46) +
      (src046[30] << 46) +
      (src046[31] << 46) +
      (src046[32] << 46) +
      (src046[33] << 46) +
      (src046[34] << 46) +
      (src046[35] << 46) +
      (src046[36] << 46) +
      (src046[37] << 46) +
      (src046[38] << 46) +
      (src046[39] << 46) +
      (src046[40] << 46) +
      (src046[41] << 46) +
      (src046[42] << 46) +
      (src046[43] << 46) +
      (src046[44] << 46) +
      (src046[45] << 46) +
      (src046[46] << 46) +
      (src047[0] << 47) +
      (src047[1] << 47) +
      (src047[2] << 47) +
      (src047[3] << 47) +
      (src047[4] << 47) +
      (src047[5] << 47) +
      (src047[6] << 47) +
      (src047[7] << 47) +
      (src047[8] << 47) +
      (src047[9] << 47) +
      (src047[10] << 47) +
      (src047[11] << 47) +
      (src047[12] << 47) +
      (src047[13] << 47) +
      (src047[14] << 47) +
      (src047[15] << 47) +
      (src047[16] << 47) +
      (src047[17] << 47) +
      (src047[18] << 47) +
      (src047[19] << 47) +
      (src047[20] << 47) +
      (src047[21] << 47) +
      (src047[22] << 47) +
      (src047[23] << 47) +
      (src047[24] << 47) +
      (src047[25] << 47) +
      (src047[26] << 47) +
      (src047[27] << 47) +
      (src047[28] << 47) +
      (src047[29] << 47) +
      (src047[30] << 47) +
      (src047[31] << 47) +
      (src047[32] << 47) +
      (src047[33] << 47) +
      (src047[34] << 47) +
      (src047[35] << 47) +
      (src047[36] << 47) +
      (src047[37] << 47) +
      (src047[38] << 47) +
      (src047[39] << 47) +
      (src047[40] << 47) +
      (src047[41] << 47) +
      (src047[42] << 47) +
      (src047[43] << 47) +
      (src047[44] << 47) +
      (src047[45] << 47) +
      (src047[46] << 47) +
      (src047[47] << 47) +
      (src048[0] << 48) +
      (src048[1] << 48) +
      (src048[2] << 48) +
      (src048[3] << 48) +
      (src048[4] << 48) +
      (src048[5] << 48) +
      (src048[6] << 48) +
      (src048[7] << 48) +
      (src048[8] << 48) +
      (src048[9] << 48) +
      (src048[10] << 48) +
      (src048[11] << 48) +
      (src048[12] << 48) +
      (src048[13] << 48) +
      (src048[14] << 48) +
      (src048[15] << 48) +
      (src048[16] << 48) +
      (src048[17] << 48) +
      (src048[18] << 48) +
      (src048[19] << 48) +
      (src048[20] << 48) +
      (src048[21] << 48) +
      (src048[22] << 48) +
      (src048[23] << 48) +
      (src048[24] << 48) +
      (src048[25] << 48) +
      (src048[26] << 48) +
      (src048[27] << 48) +
      (src048[28] << 48) +
      (src048[29] << 48) +
      (src048[30] << 48) +
      (src048[31] << 48) +
      (src048[32] << 48) +
      (src048[33] << 48) +
      (src048[34] << 48) +
      (src048[35] << 48) +
      (src048[36] << 48) +
      (src048[37] << 48) +
      (src048[38] << 48) +
      (src048[39] << 48) +
      (src048[40] << 48) +
      (src048[41] << 48) +
      (src048[42] << 48) +
      (src048[43] << 48) +
      (src048[44] << 48) +
      (src048[45] << 48) +
      (src048[46] << 48) +
      (src048[47] << 48) +
      (src048[48] << 48) +
      (src049[0] << 49) +
      (src049[1] << 49) +
      (src049[2] << 49) +
      (src049[3] << 49) +
      (src049[4] << 49) +
      (src049[5] << 49) +
      (src049[6] << 49) +
      (src049[7] << 49) +
      (src049[8] << 49) +
      (src049[9] << 49) +
      (src049[10] << 49) +
      (src049[11] << 49) +
      (src049[12] << 49) +
      (src049[13] << 49) +
      (src049[14] << 49) +
      (src049[15] << 49) +
      (src049[16] << 49) +
      (src049[17] << 49) +
      (src049[18] << 49) +
      (src049[19] << 49) +
      (src049[20] << 49) +
      (src049[21] << 49) +
      (src049[22] << 49) +
      (src049[23] << 49) +
      (src049[24] << 49) +
      (src049[25] << 49) +
      (src049[26] << 49) +
      (src049[27] << 49) +
      (src049[28] << 49) +
      (src049[29] << 49) +
      (src049[30] << 49) +
      (src049[31] << 49) +
      (src049[32] << 49) +
      (src049[33] << 49) +
      (src049[34] << 49) +
      (src049[35] << 49) +
      (src049[36] << 49) +
      (src049[37] << 49) +
      (src049[38] << 49) +
      (src049[39] << 49) +
      (src049[40] << 49) +
      (src049[41] << 49) +
      (src049[42] << 49) +
      (src049[43] << 49) +
      (src049[44] << 49) +
      (src049[45] << 49) +
      (src049[46] << 49) +
      (src049[47] << 49) +
      (src049[48] << 49) +
      (src049[49] << 49) +
      (src050[0] << 50) +
      (src050[1] << 50) +
      (src050[2] << 50) +
      (src050[3] << 50) +
      (src050[4] << 50) +
      (src050[5] << 50) +
      (src050[6] << 50) +
      (src050[7] << 50) +
      (src050[8] << 50) +
      (src050[9] << 50) +
      (src050[10] << 50) +
      (src050[11] << 50) +
      (src050[12] << 50) +
      (src050[13] << 50) +
      (src050[14] << 50) +
      (src050[15] << 50) +
      (src050[16] << 50) +
      (src050[17] << 50) +
      (src050[18] << 50) +
      (src050[19] << 50) +
      (src050[20] << 50) +
      (src050[21] << 50) +
      (src050[22] << 50) +
      (src050[23] << 50) +
      (src050[24] << 50) +
      (src050[25] << 50) +
      (src050[26] << 50) +
      (src050[27] << 50) +
      (src050[28] << 50) +
      (src050[29] << 50) +
      (src050[30] << 50) +
      (src050[31] << 50) +
      (src050[32] << 50) +
      (src050[33] << 50) +
      (src050[34] << 50) +
      (src050[35] << 50) +
      (src050[36] << 50) +
      (src050[37] << 50) +
      (src050[38] << 50) +
      (src050[39] << 50) +
      (src050[40] << 50) +
      (src050[41] << 50) +
      (src050[42] << 50) +
      (src050[43] << 50) +
      (src050[44] << 50) +
      (src050[45] << 50) +
      (src050[46] << 50) +
      (src050[47] << 50) +
      (src050[48] << 50) +
      (src050[49] << 50) +
      (src050[50] << 50) +
      (src051[0] << 51) +
      (src051[1] << 51) +
      (src051[2] << 51) +
      (src051[3] << 51) +
      (src051[4] << 51) +
      (src051[5] << 51) +
      (src051[6] << 51) +
      (src051[7] << 51) +
      (src051[8] << 51) +
      (src051[9] << 51) +
      (src051[10] << 51) +
      (src051[11] << 51) +
      (src051[12] << 51) +
      (src051[13] << 51) +
      (src051[14] << 51) +
      (src051[15] << 51) +
      (src051[16] << 51) +
      (src051[17] << 51) +
      (src051[18] << 51) +
      (src051[19] << 51) +
      (src051[20] << 51) +
      (src051[21] << 51) +
      (src051[22] << 51) +
      (src051[23] << 51) +
      (src051[24] << 51) +
      (src051[25] << 51) +
      (src051[26] << 51) +
      (src051[27] << 51) +
      (src051[28] << 51) +
      (src051[29] << 51) +
      (src051[30] << 51) +
      (src051[31] << 51) +
      (src051[32] << 51) +
      (src051[33] << 51) +
      (src051[34] << 51) +
      (src051[35] << 51) +
      (src051[36] << 51) +
      (src051[37] << 51) +
      (src051[38] << 51) +
      (src051[39] << 51) +
      (src051[40] << 51) +
      (src051[41] << 51) +
      (src051[42] << 51) +
      (src051[43] << 51) +
      (src051[44] << 51) +
      (src051[45] << 51) +
      (src051[46] << 51) +
      (src051[47] << 51) +
      (src051[48] << 51) +
      (src051[49] << 51) +
      (src051[50] << 51) +
      (src051[51] << 51) +
      (src052[0] << 52) +
      (src052[1] << 52) +
      (src052[2] << 52) +
      (src052[3] << 52) +
      (src052[4] << 52) +
      (src052[5] << 52) +
      (src052[6] << 52) +
      (src052[7] << 52) +
      (src052[8] << 52) +
      (src052[9] << 52) +
      (src052[10] << 52) +
      (src052[11] << 52) +
      (src052[12] << 52) +
      (src052[13] << 52) +
      (src052[14] << 52) +
      (src052[15] << 52) +
      (src052[16] << 52) +
      (src052[17] << 52) +
      (src052[18] << 52) +
      (src052[19] << 52) +
      (src052[20] << 52) +
      (src052[21] << 52) +
      (src052[22] << 52) +
      (src052[23] << 52) +
      (src052[24] << 52) +
      (src052[25] << 52) +
      (src052[26] << 52) +
      (src052[27] << 52) +
      (src052[28] << 52) +
      (src052[29] << 52) +
      (src052[30] << 52) +
      (src052[31] << 52) +
      (src052[32] << 52) +
      (src052[33] << 52) +
      (src052[34] << 52) +
      (src052[35] << 52) +
      (src052[36] << 52) +
      (src052[37] << 52) +
      (src052[38] << 52) +
      (src052[39] << 52) +
      (src052[40] << 52) +
      (src052[41] << 52) +
      (src052[42] << 52) +
      (src052[43] << 52) +
      (src052[44] << 52) +
      (src052[45] << 52) +
      (src052[46] << 52) +
      (src052[47] << 52) +
      (src052[48] << 52) +
      (src052[49] << 52) +
      (src052[50] << 52) +
      (src052[51] << 52) +
      (src052[52] << 52) +
      (src053[0] << 53) +
      (src053[1] << 53) +
      (src053[2] << 53) +
      (src053[3] << 53) +
      (src053[4] << 53) +
      (src053[5] << 53) +
      (src053[6] << 53) +
      (src053[7] << 53) +
      (src053[8] << 53) +
      (src053[9] << 53) +
      (src053[10] << 53) +
      (src053[11] << 53) +
      (src053[12] << 53) +
      (src053[13] << 53) +
      (src053[14] << 53) +
      (src053[15] << 53) +
      (src053[16] << 53) +
      (src053[17] << 53) +
      (src053[18] << 53) +
      (src053[19] << 53) +
      (src053[20] << 53) +
      (src053[21] << 53) +
      (src053[22] << 53) +
      (src053[23] << 53) +
      (src053[24] << 53) +
      (src053[25] << 53) +
      (src053[26] << 53) +
      (src053[27] << 53) +
      (src053[28] << 53) +
      (src053[29] << 53) +
      (src053[30] << 53) +
      (src053[31] << 53) +
      (src053[32] << 53) +
      (src053[33] << 53) +
      (src053[34] << 53) +
      (src053[35] << 53) +
      (src053[36] << 53) +
      (src053[37] << 53) +
      (src053[38] << 53) +
      (src053[39] << 53) +
      (src053[40] << 53) +
      (src053[41] << 53) +
      (src053[42] << 53) +
      (src053[43] << 53) +
      (src053[44] << 53) +
      (src053[45] << 53) +
      (src053[46] << 53) +
      (src053[47] << 53) +
      (src053[48] << 53) +
      (src053[49] << 53) +
      (src053[50] << 53) +
      (src053[51] << 53) +
      (src053[52] << 53) +
      (src053[53] << 53) +
      (src054[0] << 54) +
      (src054[1] << 54) +
      (src054[2] << 54) +
      (src054[3] << 54) +
      (src054[4] << 54) +
      (src054[5] << 54) +
      (src054[6] << 54) +
      (src054[7] << 54) +
      (src054[8] << 54) +
      (src054[9] << 54) +
      (src054[10] << 54) +
      (src054[11] << 54) +
      (src054[12] << 54) +
      (src054[13] << 54) +
      (src054[14] << 54) +
      (src054[15] << 54) +
      (src054[16] << 54) +
      (src054[17] << 54) +
      (src054[18] << 54) +
      (src054[19] << 54) +
      (src054[20] << 54) +
      (src054[21] << 54) +
      (src054[22] << 54) +
      (src054[23] << 54) +
      (src054[24] << 54) +
      (src054[25] << 54) +
      (src054[26] << 54) +
      (src054[27] << 54) +
      (src054[28] << 54) +
      (src054[29] << 54) +
      (src054[30] << 54) +
      (src054[31] << 54) +
      (src054[32] << 54) +
      (src054[33] << 54) +
      (src054[34] << 54) +
      (src054[35] << 54) +
      (src054[36] << 54) +
      (src054[37] << 54) +
      (src054[38] << 54) +
      (src054[39] << 54) +
      (src054[40] << 54) +
      (src054[41] << 54) +
      (src054[42] << 54) +
      (src054[43] << 54) +
      (src054[44] << 54) +
      (src054[45] << 54) +
      (src054[46] << 54) +
      (src054[47] << 54) +
      (src054[48] << 54) +
      (src054[49] << 54) +
      (src054[50] << 54) +
      (src054[51] << 54) +
      (src054[52] << 54) +
      (src054[53] << 54) +
      (src054[54] << 54) +
      (src055[0] << 55) +
      (src055[1] << 55) +
      (src055[2] << 55) +
      (src055[3] << 55) +
      (src055[4] << 55) +
      (src055[5] << 55) +
      (src055[6] << 55) +
      (src055[7] << 55) +
      (src055[8] << 55) +
      (src055[9] << 55) +
      (src055[10] << 55) +
      (src055[11] << 55) +
      (src055[12] << 55) +
      (src055[13] << 55) +
      (src055[14] << 55) +
      (src055[15] << 55) +
      (src055[16] << 55) +
      (src055[17] << 55) +
      (src055[18] << 55) +
      (src055[19] << 55) +
      (src055[20] << 55) +
      (src055[21] << 55) +
      (src055[22] << 55) +
      (src055[23] << 55) +
      (src055[24] << 55) +
      (src055[25] << 55) +
      (src055[26] << 55) +
      (src055[27] << 55) +
      (src055[28] << 55) +
      (src055[29] << 55) +
      (src055[30] << 55) +
      (src055[31] << 55) +
      (src055[32] << 55) +
      (src055[33] << 55) +
      (src055[34] << 55) +
      (src055[35] << 55) +
      (src055[36] << 55) +
      (src055[37] << 55) +
      (src055[38] << 55) +
      (src055[39] << 55) +
      (src055[40] << 55) +
      (src055[41] << 55) +
      (src055[42] << 55) +
      (src055[43] << 55) +
      (src055[44] << 55) +
      (src055[45] << 55) +
      (src055[46] << 55) +
      (src055[47] << 55) +
      (src055[48] << 55) +
      (src055[49] << 55) +
      (src055[50] << 55) +
      (src055[51] << 55) +
      (src055[52] << 55) +
      (src055[53] << 55) +
      (src055[54] << 55) +
      (src055[55] << 55) +
      (src056[0] << 56) +
      (src056[1] << 56) +
      (src056[2] << 56) +
      (src056[3] << 56) +
      (src056[4] << 56) +
      (src056[5] << 56) +
      (src056[6] << 56) +
      (src056[7] << 56) +
      (src056[8] << 56) +
      (src056[9] << 56) +
      (src056[10] << 56) +
      (src056[11] << 56) +
      (src056[12] << 56) +
      (src056[13] << 56) +
      (src056[14] << 56) +
      (src056[15] << 56) +
      (src056[16] << 56) +
      (src056[17] << 56) +
      (src056[18] << 56) +
      (src056[19] << 56) +
      (src056[20] << 56) +
      (src056[21] << 56) +
      (src056[22] << 56) +
      (src056[23] << 56) +
      (src056[24] << 56) +
      (src056[25] << 56) +
      (src056[26] << 56) +
      (src056[27] << 56) +
      (src056[28] << 56) +
      (src056[29] << 56) +
      (src056[30] << 56) +
      (src056[31] << 56) +
      (src056[32] << 56) +
      (src056[33] << 56) +
      (src056[34] << 56) +
      (src056[35] << 56) +
      (src056[36] << 56) +
      (src056[37] << 56) +
      (src056[38] << 56) +
      (src056[39] << 56) +
      (src056[40] << 56) +
      (src056[41] << 56) +
      (src056[42] << 56) +
      (src056[43] << 56) +
      (src056[44] << 56) +
      (src056[45] << 56) +
      (src056[46] << 56) +
      (src056[47] << 56) +
      (src056[48] << 56) +
      (src056[49] << 56) +
      (src056[50] << 56) +
      (src056[51] << 56) +
      (src056[52] << 56) +
      (src056[53] << 56) +
      (src056[54] << 56) +
      (src056[55] << 56) +
      (src056[56] << 56) +
      (src057[0] << 57) +
      (src057[1] << 57) +
      (src057[2] << 57) +
      (src057[3] << 57) +
      (src057[4] << 57) +
      (src057[5] << 57) +
      (src057[6] << 57) +
      (src057[7] << 57) +
      (src057[8] << 57) +
      (src057[9] << 57) +
      (src057[10] << 57) +
      (src057[11] << 57) +
      (src057[12] << 57) +
      (src057[13] << 57) +
      (src057[14] << 57) +
      (src057[15] << 57) +
      (src057[16] << 57) +
      (src057[17] << 57) +
      (src057[18] << 57) +
      (src057[19] << 57) +
      (src057[20] << 57) +
      (src057[21] << 57) +
      (src057[22] << 57) +
      (src057[23] << 57) +
      (src057[24] << 57) +
      (src057[25] << 57) +
      (src057[26] << 57) +
      (src057[27] << 57) +
      (src057[28] << 57) +
      (src057[29] << 57) +
      (src057[30] << 57) +
      (src057[31] << 57) +
      (src057[32] << 57) +
      (src057[33] << 57) +
      (src057[34] << 57) +
      (src057[35] << 57) +
      (src057[36] << 57) +
      (src057[37] << 57) +
      (src057[38] << 57) +
      (src057[39] << 57) +
      (src057[40] << 57) +
      (src057[41] << 57) +
      (src057[42] << 57) +
      (src057[43] << 57) +
      (src057[44] << 57) +
      (src057[45] << 57) +
      (src057[46] << 57) +
      (src057[47] << 57) +
      (src057[48] << 57) +
      (src057[49] << 57) +
      (src057[50] << 57) +
      (src057[51] << 57) +
      (src057[52] << 57) +
      (src057[53] << 57) +
      (src057[54] << 57) +
      (src057[55] << 57) +
      (src057[56] << 57) +
      (src057[57] << 57) +
      (src058[0] << 58) +
      (src058[1] << 58) +
      (src058[2] << 58) +
      (src058[3] << 58) +
      (src058[4] << 58) +
      (src058[5] << 58) +
      (src058[6] << 58) +
      (src058[7] << 58) +
      (src058[8] << 58) +
      (src058[9] << 58) +
      (src058[10] << 58) +
      (src058[11] << 58) +
      (src058[12] << 58) +
      (src058[13] << 58) +
      (src058[14] << 58) +
      (src058[15] << 58) +
      (src058[16] << 58) +
      (src058[17] << 58) +
      (src058[18] << 58) +
      (src058[19] << 58) +
      (src058[20] << 58) +
      (src058[21] << 58) +
      (src058[22] << 58) +
      (src058[23] << 58) +
      (src058[24] << 58) +
      (src058[25] << 58) +
      (src058[26] << 58) +
      (src058[27] << 58) +
      (src058[28] << 58) +
      (src058[29] << 58) +
      (src058[30] << 58) +
      (src058[31] << 58) +
      (src058[32] << 58) +
      (src058[33] << 58) +
      (src058[34] << 58) +
      (src058[35] << 58) +
      (src058[36] << 58) +
      (src058[37] << 58) +
      (src058[38] << 58) +
      (src058[39] << 58) +
      (src058[40] << 58) +
      (src058[41] << 58) +
      (src058[42] << 58) +
      (src058[43] << 58) +
      (src058[44] << 58) +
      (src058[45] << 58) +
      (src058[46] << 58) +
      (src058[47] << 58) +
      (src058[48] << 58) +
      (src058[49] << 58) +
      (src058[50] << 58) +
      (src058[51] << 58) +
      (src058[52] << 58) +
      (src058[53] << 58) +
      (src058[54] << 58) +
      (src058[55] << 58) +
      (src058[56] << 58) +
      (src058[57] << 58) +
      (src058[58] << 58) +
      (src059[0] << 59) +
      (src059[1] << 59) +
      (src059[2] << 59) +
      (src059[3] << 59) +
      (src059[4] << 59) +
      (src059[5] << 59) +
      (src059[6] << 59) +
      (src059[7] << 59) +
      (src059[8] << 59) +
      (src059[9] << 59) +
      (src059[10] << 59) +
      (src059[11] << 59) +
      (src059[12] << 59) +
      (src059[13] << 59) +
      (src059[14] << 59) +
      (src059[15] << 59) +
      (src059[16] << 59) +
      (src059[17] << 59) +
      (src059[18] << 59) +
      (src059[19] << 59) +
      (src059[20] << 59) +
      (src059[21] << 59) +
      (src059[22] << 59) +
      (src059[23] << 59) +
      (src059[24] << 59) +
      (src059[25] << 59) +
      (src059[26] << 59) +
      (src059[27] << 59) +
      (src059[28] << 59) +
      (src059[29] << 59) +
      (src059[30] << 59) +
      (src059[31] << 59) +
      (src059[32] << 59) +
      (src059[33] << 59) +
      (src059[34] << 59) +
      (src059[35] << 59) +
      (src059[36] << 59) +
      (src059[37] << 59) +
      (src059[38] << 59) +
      (src059[39] << 59) +
      (src059[40] << 59) +
      (src059[41] << 59) +
      (src059[42] << 59) +
      (src059[43] << 59) +
      (src059[44] << 59) +
      (src059[45] << 59) +
      (src059[46] << 59) +
      (src059[47] << 59) +
      (src059[48] << 59) +
      (src059[49] << 59) +
      (src059[50] << 59) +
      (src059[51] << 59) +
      (src059[52] << 59) +
      (src059[53] << 59) +
      (src059[54] << 59) +
      (src059[55] << 59) +
      (src059[56] << 59) +
      (src059[57] << 59) +
      (src059[58] << 59) +
      (src059[59] << 59) +
      (src060[0] << 60) +
      (src060[1] << 60) +
      (src060[2] << 60) +
      (src060[3] << 60) +
      (src060[4] << 60) +
      (src060[5] << 60) +
      (src060[6] << 60) +
      (src060[7] << 60) +
      (src060[8] << 60) +
      (src060[9] << 60) +
      (src060[10] << 60) +
      (src060[11] << 60) +
      (src060[12] << 60) +
      (src060[13] << 60) +
      (src060[14] << 60) +
      (src060[15] << 60) +
      (src060[16] << 60) +
      (src060[17] << 60) +
      (src060[18] << 60) +
      (src060[19] << 60) +
      (src060[20] << 60) +
      (src060[21] << 60) +
      (src060[22] << 60) +
      (src060[23] << 60) +
      (src060[24] << 60) +
      (src060[25] << 60) +
      (src060[26] << 60) +
      (src060[27] << 60) +
      (src060[28] << 60) +
      (src060[29] << 60) +
      (src060[30] << 60) +
      (src060[31] << 60) +
      (src060[32] << 60) +
      (src060[33] << 60) +
      (src060[34] << 60) +
      (src060[35] << 60) +
      (src060[36] << 60) +
      (src060[37] << 60) +
      (src060[38] << 60) +
      (src060[39] << 60) +
      (src060[40] << 60) +
      (src060[41] << 60) +
      (src060[42] << 60) +
      (src060[43] << 60) +
      (src060[44] << 60) +
      (src060[45] << 60) +
      (src060[46] << 60) +
      (src060[47] << 60) +
      (src060[48] << 60) +
      (src060[49] << 60) +
      (src060[50] << 60) +
      (src060[51] << 60) +
      (src060[52] << 60) +
      (src060[53] << 60) +
      (src060[54] << 60) +
      (src060[55] << 60) +
      (src060[56] << 60) +
      (src060[57] << 60) +
      (src060[58] << 60) +
      (src060[59] << 60) +
      (src060[60] << 60) +
      (src061[0] << 61) +
      (src061[1] << 61) +
      (src061[2] << 61) +
      (src061[3] << 61) +
      (src061[4] << 61) +
      (src061[5] << 61) +
      (src061[6] << 61) +
      (src061[7] << 61) +
      (src061[8] << 61) +
      (src061[9] << 61) +
      (src061[10] << 61) +
      (src061[11] << 61) +
      (src061[12] << 61) +
      (src061[13] << 61) +
      (src061[14] << 61) +
      (src061[15] << 61) +
      (src061[16] << 61) +
      (src061[17] << 61) +
      (src061[18] << 61) +
      (src061[19] << 61) +
      (src061[20] << 61) +
      (src061[21] << 61) +
      (src061[22] << 61) +
      (src061[23] << 61) +
      (src061[24] << 61) +
      (src061[25] << 61) +
      (src061[26] << 61) +
      (src061[27] << 61) +
      (src061[28] << 61) +
      (src061[29] << 61) +
      (src061[30] << 61) +
      (src061[31] << 61) +
      (src061[32] << 61) +
      (src061[33] << 61) +
      (src061[34] << 61) +
      (src061[35] << 61) +
      (src061[36] << 61) +
      (src061[37] << 61) +
      (src061[38] << 61) +
      (src061[39] << 61) +
      (src061[40] << 61) +
      (src061[41] << 61) +
      (src061[42] << 61) +
      (src061[43] << 61) +
      (src061[44] << 61) +
      (src061[45] << 61) +
      (src061[46] << 61) +
      (src061[47] << 61) +
      (src061[48] << 61) +
      (src061[49] << 61) +
      (src061[50] << 61) +
      (src061[51] << 61) +
      (src061[52] << 61) +
      (src061[53] << 61) +
      (src061[54] << 61) +
      (src061[55] << 61) +
      (src061[56] << 61) +
      (src061[57] << 61) +
      (src061[58] << 61) +
      (src061[59] << 61) +
      (src061[60] << 61) +
      (src061[61] << 61) +
      (src062[0] << 62) +
      (src062[1] << 62) +
      (src062[2] << 62) +
      (src062[3] << 62) +
      (src062[4] << 62) +
      (src062[5] << 62) +
      (src062[6] << 62) +
      (src062[7] << 62) +
      (src062[8] << 62) +
      (src062[9] << 62) +
      (src062[10] << 62) +
      (src062[11] << 62) +
      (src062[12] << 62) +
      (src062[13] << 62) +
      (src062[14] << 62) +
      (src062[15] << 62) +
      (src062[16] << 62) +
      (src062[17] << 62) +
      (src062[18] << 62) +
      (src062[19] << 62) +
      (src062[20] << 62) +
      (src062[21] << 62) +
      (src062[22] << 62) +
      (src062[23] << 62) +
      (src062[24] << 62) +
      (src062[25] << 62) +
      (src062[26] << 62) +
      (src062[27] << 62) +
      (src062[28] << 62) +
      (src062[29] << 62) +
      (src062[30] << 62) +
      (src062[31] << 62) +
      (src062[32] << 62) +
      (src062[33] << 62) +
      (src062[34] << 62) +
      (src062[35] << 62) +
      (src062[36] << 62) +
      (src062[37] << 62) +
      (src062[38] << 62) +
      (src062[39] << 62) +
      (src062[40] << 62) +
      (src062[41] << 62) +
      (src062[42] << 62) +
      (src062[43] << 62) +
      (src062[44] << 62) +
      (src062[45] << 62) +
      (src062[46] << 62) +
      (src062[47] << 62) +
      (src062[48] << 62) +
      (src062[49] << 62) +
      (src062[50] << 62) +
      (src062[51] << 62) +
      (src062[52] << 62) +
      (src062[53] << 62) +
      (src062[54] << 62) +
      (src062[55] << 62) +
      (src062[56] << 62) +
      (src062[57] << 62) +
      (src062[58] << 62) +
      (src062[59] << 62) +
      (src062[60] << 62) +
      (src062[61] << 62) +
      (src062[62] << 62) +
      (src063[0] << 63) +
      (src063[1] << 63) +
      (src063[2] << 63) +
      (src063[3] << 63) +
      (src063[4] << 63) +
      (src063[5] << 63) +
      (src063[6] << 63) +
      (src063[7] << 63) +
      (src063[8] << 63) +
      (src063[9] << 63) +
      (src063[10] << 63) +
      (src063[11] << 63) +
      (src063[12] << 63) +
      (src063[13] << 63) +
      (src063[14] << 63) +
      (src063[15] << 63) +
      (src063[16] << 63) +
      (src063[17] << 63) +
      (src063[18] << 63) +
      (src063[19] << 63) +
      (src063[20] << 63) +
      (src063[21] << 63) +
      (src063[22] << 63) +
      (src063[23] << 63) +
      (src063[24] << 63) +
      (src063[25] << 63) +
      (src063[26] << 63) +
      (src063[27] << 63) +
      (src063[28] << 63) +
      (src063[29] << 63) +
      (src063[30] << 63) +
      (src063[31] << 63) +
      (src063[32] << 63) +
      (src063[33] << 63) +
      (src063[34] << 63) +
      (src063[35] << 63) +
      (src063[36] << 63) +
      (src063[37] << 63) +
      (src063[38] << 63) +
      (src063[39] << 63) +
      (src063[40] << 63) +
      (src063[41] << 63) +
      (src063[42] << 63) +
      (src063[43] << 63) +
      (src063[44] << 63) +
      (src063[45] << 63) +
      (src063[46] << 63) +
      (src063[47] << 63) +
      (src063[48] << 63) +
      (src063[49] << 63) +
      (src063[50] << 63) +
      (src063[51] << 63) +
      (src063[52] << 63) +
      (src063[53] << 63) +
      (src063[54] << 63) +
      (src063[55] << 63) +
      (src063[56] << 63) +
      (src063[57] << 63) +
      (src063[58] << 63) +
      (src063[59] << 63) +
      (src063[60] << 63) +
      (src063[61] << 63) +
      (src063[62] << 63) +
      (src063[63] << 63) +
      (src064[0] << 64) +
      (src064[1] << 64) +
      (src064[2] << 64) +
      (src064[3] << 64) +
      (src064[4] << 64) +
      (src064[5] << 64) +
      (src064[6] << 64) +
      (src064[7] << 64) +
      (src064[8] << 64) +
      (src064[9] << 64) +
      (src064[10] << 64) +
      (src064[11] << 64) +
      (src064[12] << 64) +
      (src064[13] << 64) +
      (src064[14] << 64) +
      (src064[15] << 64) +
      (src064[16] << 64) +
      (src064[17] << 64) +
      (src064[18] << 64) +
      (src064[19] << 64) +
      (src064[20] << 64) +
      (src064[21] << 64) +
      (src064[22] << 64) +
      (src064[23] << 64) +
      (src064[24] << 64) +
      (src064[25] << 64) +
      (src064[26] << 64) +
      (src064[27] << 64) +
      (src064[28] << 64) +
      (src064[29] << 64) +
      (src064[30] << 64) +
      (src064[31] << 64) +
      (src064[32] << 64) +
      (src064[33] << 64) +
      (src064[34] << 64) +
      (src064[35] << 64) +
      (src064[36] << 64) +
      (src064[37] << 64) +
      (src064[38] << 64) +
      (src064[39] << 64) +
      (src064[40] << 64) +
      (src064[41] << 64) +
      (src064[42] << 64) +
      (src064[43] << 64) +
      (src064[44] << 64) +
      (src064[45] << 64) +
      (src064[46] << 64) +
      (src064[47] << 64) +
      (src064[48] << 64) +
      (src064[49] << 64) +
      (src064[50] << 64) +
      (src064[51] << 64) +
      (src064[52] << 64) +
      (src064[53] << 64) +
      (src064[54] << 64) +
      (src064[55] << 64) +
      (src064[56] << 64) +
      (src064[57] << 64) +
      (src064[58] << 64) +
      (src064[59] << 64) +
      (src064[60] << 64) +
      (src064[61] << 64) +
      (src064[62] << 64) +
      (src065[0] << 65) +
      (src065[1] << 65) +
      (src065[2] << 65) +
      (src065[3] << 65) +
      (src065[4] << 65) +
      (src065[5] << 65) +
      (src065[6] << 65) +
      (src065[7] << 65) +
      (src065[8] << 65) +
      (src065[9] << 65) +
      (src065[10] << 65) +
      (src065[11] << 65) +
      (src065[12] << 65) +
      (src065[13] << 65) +
      (src065[14] << 65) +
      (src065[15] << 65) +
      (src065[16] << 65) +
      (src065[17] << 65) +
      (src065[18] << 65) +
      (src065[19] << 65) +
      (src065[20] << 65) +
      (src065[21] << 65) +
      (src065[22] << 65) +
      (src065[23] << 65) +
      (src065[24] << 65) +
      (src065[25] << 65) +
      (src065[26] << 65) +
      (src065[27] << 65) +
      (src065[28] << 65) +
      (src065[29] << 65) +
      (src065[30] << 65) +
      (src065[31] << 65) +
      (src065[32] << 65) +
      (src065[33] << 65) +
      (src065[34] << 65) +
      (src065[35] << 65) +
      (src065[36] << 65) +
      (src065[37] << 65) +
      (src065[38] << 65) +
      (src065[39] << 65) +
      (src065[40] << 65) +
      (src065[41] << 65) +
      (src065[42] << 65) +
      (src065[43] << 65) +
      (src065[44] << 65) +
      (src065[45] << 65) +
      (src065[46] << 65) +
      (src065[47] << 65) +
      (src065[48] << 65) +
      (src065[49] << 65) +
      (src065[50] << 65) +
      (src065[51] << 65) +
      (src065[52] << 65) +
      (src065[53] << 65) +
      (src065[54] << 65) +
      (src065[55] << 65) +
      (src065[56] << 65) +
      (src065[57] << 65) +
      (src065[58] << 65) +
      (src065[59] << 65) +
      (src065[60] << 65) +
      (src065[61] << 65) +
      (src066[0] << 66) +
      (src066[1] << 66) +
      (src066[2] << 66) +
      (src066[3] << 66) +
      (src066[4] << 66) +
      (src066[5] << 66) +
      (src066[6] << 66) +
      (src066[7] << 66) +
      (src066[8] << 66) +
      (src066[9] << 66) +
      (src066[10] << 66) +
      (src066[11] << 66) +
      (src066[12] << 66) +
      (src066[13] << 66) +
      (src066[14] << 66) +
      (src066[15] << 66) +
      (src066[16] << 66) +
      (src066[17] << 66) +
      (src066[18] << 66) +
      (src066[19] << 66) +
      (src066[20] << 66) +
      (src066[21] << 66) +
      (src066[22] << 66) +
      (src066[23] << 66) +
      (src066[24] << 66) +
      (src066[25] << 66) +
      (src066[26] << 66) +
      (src066[27] << 66) +
      (src066[28] << 66) +
      (src066[29] << 66) +
      (src066[30] << 66) +
      (src066[31] << 66) +
      (src066[32] << 66) +
      (src066[33] << 66) +
      (src066[34] << 66) +
      (src066[35] << 66) +
      (src066[36] << 66) +
      (src066[37] << 66) +
      (src066[38] << 66) +
      (src066[39] << 66) +
      (src066[40] << 66) +
      (src066[41] << 66) +
      (src066[42] << 66) +
      (src066[43] << 66) +
      (src066[44] << 66) +
      (src066[45] << 66) +
      (src066[46] << 66) +
      (src066[47] << 66) +
      (src066[48] << 66) +
      (src066[49] << 66) +
      (src066[50] << 66) +
      (src066[51] << 66) +
      (src066[52] << 66) +
      (src066[53] << 66) +
      (src066[54] << 66) +
      (src066[55] << 66) +
      (src066[56] << 66) +
      (src066[57] << 66) +
      (src066[58] << 66) +
      (src066[59] << 66) +
      (src066[60] << 66) +
      (src067[0] << 67) +
      (src067[1] << 67) +
      (src067[2] << 67) +
      (src067[3] << 67) +
      (src067[4] << 67) +
      (src067[5] << 67) +
      (src067[6] << 67) +
      (src067[7] << 67) +
      (src067[8] << 67) +
      (src067[9] << 67) +
      (src067[10] << 67) +
      (src067[11] << 67) +
      (src067[12] << 67) +
      (src067[13] << 67) +
      (src067[14] << 67) +
      (src067[15] << 67) +
      (src067[16] << 67) +
      (src067[17] << 67) +
      (src067[18] << 67) +
      (src067[19] << 67) +
      (src067[20] << 67) +
      (src067[21] << 67) +
      (src067[22] << 67) +
      (src067[23] << 67) +
      (src067[24] << 67) +
      (src067[25] << 67) +
      (src067[26] << 67) +
      (src067[27] << 67) +
      (src067[28] << 67) +
      (src067[29] << 67) +
      (src067[30] << 67) +
      (src067[31] << 67) +
      (src067[32] << 67) +
      (src067[33] << 67) +
      (src067[34] << 67) +
      (src067[35] << 67) +
      (src067[36] << 67) +
      (src067[37] << 67) +
      (src067[38] << 67) +
      (src067[39] << 67) +
      (src067[40] << 67) +
      (src067[41] << 67) +
      (src067[42] << 67) +
      (src067[43] << 67) +
      (src067[44] << 67) +
      (src067[45] << 67) +
      (src067[46] << 67) +
      (src067[47] << 67) +
      (src067[48] << 67) +
      (src067[49] << 67) +
      (src067[50] << 67) +
      (src067[51] << 67) +
      (src067[52] << 67) +
      (src067[53] << 67) +
      (src067[54] << 67) +
      (src067[55] << 67) +
      (src067[56] << 67) +
      (src067[57] << 67) +
      (src067[58] << 67) +
      (src067[59] << 67) +
      (src068[0] << 68) +
      (src068[1] << 68) +
      (src068[2] << 68) +
      (src068[3] << 68) +
      (src068[4] << 68) +
      (src068[5] << 68) +
      (src068[6] << 68) +
      (src068[7] << 68) +
      (src068[8] << 68) +
      (src068[9] << 68) +
      (src068[10] << 68) +
      (src068[11] << 68) +
      (src068[12] << 68) +
      (src068[13] << 68) +
      (src068[14] << 68) +
      (src068[15] << 68) +
      (src068[16] << 68) +
      (src068[17] << 68) +
      (src068[18] << 68) +
      (src068[19] << 68) +
      (src068[20] << 68) +
      (src068[21] << 68) +
      (src068[22] << 68) +
      (src068[23] << 68) +
      (src068[24] << 68) +
      (src068[25] << 68) +
      (src068[26] << 68) +
      (src068[27] << 68) +
      (src068[28] << 68) +
      (src068[29] << 68) +
      (src068[30] << 68) +
      (src068[31] << 68) +
      (src068[32] << 68) +
      (src068[33] << 68) +
      (src068[34] << 68) +
      (src068[35] << 68) +
      (src068[36] << 68) +
      (src068[37] << 68) +
      (src068[38] << 68) +
      (src068[39] << 68) +
      (src068[40] << 68) +
      (src068[41] << 68) +
      (src068[42] << 68) +
      (src068[43] << 68) +
      (src068[44] << 68) +
      (src068[45] << 68) +
      (src068[46] << 68) +
      (src068[47] << 68) +
      (src068[48] << 68) +
      (src068[49] << 68) +
      (src068[50] << 68) +
      (src068[51] << 68) +
      (src068[52] << 68) +
      (src068[53] << 68) +
      (src068[54] << 68) +
      (src068[55] << 68) +
      (src068[56] << 68) +
      (src068[57] << 68) +
      (src068[58] << 68) +
      (src069[0] << 69) +
      (src069[1] << 69) +
      (src069[2] << 69) +
      (src069[3] << 69) +
      (src069[4] << 69) +
      (src069[5] << 69) +
      (src069[6] << 69) +
      (src069[7] << 69) +
      (src069[8] << 69) +
      (src069[9] << 69) +
      (src069[10] << 69) +
      (src069[11] << 69) +
      (src069[12] << 69) +
      (src069[13] << 69) +
      (src069[14] << 69) +
      (src069[15] << 69) +
      (src069[16] << 69) +
      (src069[17] << 69) +
      (src069[18] << 69) +
      (src069[19] << 69) +
      (src069[20] << 69) +
      (src069[21] << 69) +
      (src069[22] << 69) +
      (src069[23] << 69) +
      (src069[24] << 69) +
      (src069[25] << 69) +
      (src069[26] << 69) +
      (src069[27] << 69) +
      (src069[28] << 69) +
      (src069[29] << 69) +
      (src069[30] << 69) +
      (src069[31] << 69) +
      (src069[32] << 69) +
      (src069[33] << 69) +
      (src069[34] << 69) +
      (src069[35] << 69) +
      (src069[36] << 69) +
      (src069[37] << 69) +
      (src069[38] << 69) +
      (src069[39] << 69) +
      (src069[40] << 69) +
      (src069[41] << 69) +
      (src069[42] << 69) +
      (src069[43] << 69) +
      (src069[44] << 69) +
      (src069[45] << 69) +
      (src069[46] << 69) +
      (src069[47] << 69) +
      (src069[48] << 69) +
      (src069[49] << 69) +
      (src069[50] << 69) +
      (src069[51] << 69) +
      (src069[52] << 69) +
      (src069[53] << 69) +
      (src069[54] << 69) +
      (src069[55] << 69) +
      (src069[56] << 69) +
      (src069[57] << 69) +
      (src070[0] << 70) +
      (src070[1] << 70) +
      (src070[2] << 70) +
      (src070[3] << 70) +
      (src070[4] << 70) +
      (src070[5] << 70) +
      (src070[6] << 70) +
      (src070[7] << 70) +
      (src070[8] << 70) +
      (src070[9] << 70) +
      (src070[10] << 70) +
      (src070[11] << 70) +
      (src070[12] << 70) +
      (src070[13] << 70) +
      (src070[14] << 70) +
      (src070[15] << 70) +
      (src070[16] << 70) +
      (src070[17] << 70) +
      (src070[18] << 70) +
      (src070[19] << 70) +
      (src070[20] << 70) +
      (src070[21] << 70) +
      (src070[22] << 70) +
      (src070[23] << 70) +
      (src070[24] << 70) +
      (src070[25] << 70) +
      (src070[26] << 70) +
      (src070[27] << 70) +
      (src070[28] << 70) +
      (src070[29] << 70) +
      (src070[30] << 70) +
      (src070[31] << 70) +
      (src070[32] << 70) +
      (src070[33] << 70) +
      (src070[34] << 70) +
      (src070[35] << 70) +
      (src070[36] << 70) +
      (src070[37] << 70) +
      (src070[38] << 70) +
      (src070[39] << 70) +
      (src070[40] << 70) +
      (src070[41] << 70) +
      (src070[42] << 70) +
      (src070[43] << 70) +
      (src070[44] << 70) +
      (src070[45] << 70) +
      (src070[46] << 70) +
      (src070[47] << 70) +
      (src070[48] << 70) +
      (src070[49] << 70) +
      (src070[50] << 70) +
      (src070[51] << 70) +
      (src070[52] << 70) +
      (src070[53] << 70) +
      (src070[54] << 70) +
      (src070[55] << 70) +
      (src070[56] << 70) +
      (src071[0] << 71) +
      (src071[1] << 71) +
      (src071[2] << 71) +
      (src071[3] << 71) +
      (src071[4] << 71) +
      (src071[5] << 71) +
      (src071[6] << 71) +
      (src071[7] << 71) +
      (src071[8] << 71) +
      (src071[9] << 71) +
      (src071[10] << 71) +
      (src071[11] << 71) +
      (src071[12] << 71) +
      (src071[13] << 71) +
      (src071[14] << 71) +
      (src071[15] << 71) +
      (src071[16] << 71) +
      (src071[17] << 71) +
      (src071[18] << 71) +
      (src071[19] << 71) +
      (src071[20] << 71) +
      (src071[21] << 71) +
      (src071[22] << 71) +
      (src071[23] << 71) +
      (src071[24] << 71) +
      (src071[25] << 71) +
      (src071[26] << 71) +
      (src071[27] << 71) +
      (src071[28] << 71) +
      (src071[29] << 71) +
      (src071[30] << 71) +
      (src071[31] << 71) +
      (src071[32] << 71) +
      (src071[33] << 71) +
      (src071[34] << 71) +
      (src071[35] << 71) +
      (src071[36] << 71) +
      (src071[37] << 71) +
      (src071[38] << 71) +
      (src071[39] << 71) +
      (src071[40] << 71) +
      (src071[41] << 71) +
      (src071[42] << 71) +
      (src071[43] << 71) +
      (src071[44] << 71) +
      (src071[45] << 71) +
      (src071[46] << 71) +
      (src071[47] << 71) +
      (src071[48] << 71) +
      (src071[49] << 71) +
      (src071[50] << 71) +
      (src071[51] << 71) +
      (src071[52] << 71) +
      (src071[53] << 71) +
      (src071[54] << 71) +
      (src071[55] << 71) +
      (src072[0] << 72) +
      (src072[1] << 72) +
      (src072[2] << 72) +
      (src072[3] << 72) +
      (src072[4] << 72) +
      (src072[5] << 72) +
      (src072[6] << 72) +
      (src072[7] << 72) +
      (src072[8] << 72) +
      (src072[9] << 72) +
      (src072[10] << 72) +
      (src072[11] << 72) +
      (src072[12] << 72) +
      (src072[13] << 72) +
      (src072[14] << 72) +
      (src072[15] << 72) +
      (src072[16] << 72) +
      (src072[17] << 72) +
      (src072[18] << 72) +
      (src072[19] << 72) +
      (src072[20] << 72) +
      (src072[21] << 72) +
      (src072[22] << 72) +
      (src072[23] << 72) +
      (src072[24] << 72) +
      (src072[25] << 72) +
      (src072[26] << 72) +
      (src072[27] << 72) +
      (src072[28] << 72) +
      (src072[29] << 72) +
      (src072[30] << 72) +
      (src072[31] << 72) +
      (src072[32] << 72) +
      (src072[33] << 72) +
      (src072[34] << 72) +
      (src072[35] << 72) +
      (src072[36] << 72) +
      (src072[37] << 72) +
      (src072[38] << 72) +
      (src072[39] << 72) +
      (src072[40] << 72) +
      (src072[41] << 72) +
      (src072[42] << 72) +
      (src072[43] << 72) +
      (src072[44] << 72) +
      (src072[45] << 72) +
      (src072[46] << 72) +
      (src072[47] << 72) +
      (src072[48] << 72) +
      (src072[49] << 72) +
      (src072[50] << 72) +
      (src072[51] << 72) +
      (src072[52] << 72) +
      (src072[53] << 72) +
      (src072[54] << 72) +
      (src073[0] << 73) +
      (src073[1] << 73) +
      (src073[2] << 73) +
      (src073[3] << 73) +
      (src073[4] << 73) +
      (src073[5] << 73) +
      (src073[6] << 73) +
      (src073[7] << 73) +
      (src073[8] << 73) +
      (src073[9] << 73) +
      (src073[10] << 73) +
      (src073[11] << 73) +
      (src073[12] << 73) +
      (src073[13] << 73) +
      (src073[14] << 73) +
      (src073[15] << 73) +
      (src073[16] << 73) +
      (src073[17] << 73) +
      (src073[18] << 73) +
      (src073[19] << 73) +
      (src073[20] << 73) +
      (src073[21] << 73) +
      (src073[22] << 73) +
      (src073[23] << 73) +
      (src073[24] << 73) +
      (src073[25] << 73) +
      (src073[26] << 73) +
      (src073[27] << 73) +
      (src073[28] << 73) +
      (src073[29] << 73) +
      (src073[30] << 73) +
      (src073[31] << 73) +
      (src073[32] << 73) +
      (src073[33] << 73) +
      (src073[34] << 73) +
      (src073[35] << 73) +
      (src073[36] << 73) +
      (src073[37] << 73) +
      (src073[38] << 73) +
      (src073[39] << 73) +
      (src073[40] << 73) +
      (src073[41] << 73) +
      (src073[42] << 73) +
      (src073[43] << 73) +
      (src073[44] << 73) +
      (src073[45] << 73) +
      (src073[46] << 73) +
      (src073[47] << 73) +
      (src073[48] << 73) +
      (src073[49] << 73) +
      (src073[50] << 73) +
      (src073[51] << 73) +
      (src073[52] << 73) +
      (src073[53] << 73) +
      (src074[0] << 74) +
      (src074[1] << 74) +
      (src074[2] << 74) +
      (src074[3] << 74) +
      (src074[4] << 74) +
      (src074[5] << 74) +
      (src074[6] << 74) +
      (src074[7] << 74) +
      (src074[8] << 74) +
      (src074[9] << 74) +
      (src074[10] << 74) +
      (src074[11] << 74) +
      (src074[12] << 74) +
      (src074[13] << 74) +
      (src074[14] << 74) +
      (src074[15] << 74) +
      (src074[16] << 74) +
      (src074[17] << 74) +
      (src074[18] << 74) +
      (src074[19] << 74) +
      (src074[20] << 74) +
      (src074[21] << 74) +
      (src074[22] << 74) +
      (src074[23] << 74) +
      (src074[24] << 74) +
      (src074[25] << 74) +
      (src074[26] << 74) +
      (src074[27] << 74) +
      (src074[28] << 74) +
      (src074[29] << 74) +
      (src074[30] << 74) +
      (src074[31] << 74) +
      (src074[32] << 74) +
      (src074[33] << 74) +
      (src074[34] << 74) +
      (src074[35] << 74) +
      (src074[36] << 74) +
      (src074[37] << 74) +
      (src074[38] << 74) +
      (src074[39] << 74) +
      (src074[40] << 74) +
      (src074[41] << 74) +
      (src074[42] << 74) +
      (src074[43] << 74) +
      (src074[44] << 74) +
      (src074[45] << 74) +
      (src074[46] << 74) +
      (src074[47] << 74) +
      (src074[48] << 74) +
      (src074[49] << 74) +
      (src074[50] << 74) +
      (src074[51] << 74) +
      (src074[52] << 74) +
      (src075[0] << 75) +
      (src075[1] << 75) +
      (src075[2] << 75) +
      (src075[3] << 75) +
      (src075[4] << 75) +
      (src075[5] << 75) +
      (src075[6] << 75) +
      (src075[7] << 75) +
      (src075[8] << 75) +
      (src075[9] << 75) +
      (src075[10] << 75) +
      (src075[11] << 75) +
      (src075[12] << 75) +
      (src075[13] << 75) +
      (src075[14] << 75) +
      (src075[15] << 75) +
      (src075[16] << 75) +
      (src075[17] << 75) +
      (src075[18] << 75) +
      (src075[19] << 75) +
      (src075[20] << 75) +
      (src075[21] << 75) +
      (src075[22] << 75) +
      (src075[23] << 75) +
      (src075[24] << 75) +
      (src075[25] << 75) +
      (src075[26] << 75) +
      (src075[27] << 75) +
      (src075[28] << 75) +
      (src075[29] << 75) +
      (src075[30] << 75) +
      (src075[31] << 75) +
      (src075[32] << 75) +
      (src075[33] << 75) +
      (src075[34] << 75) +
      (src075[35] << 75) +
      (src075[36] << 75) +
      (src075[37] << 75) +
      (src075[38] << 75) +
      (src075[39] << 75) +
      (src075[40] << 75) +
      (src075[41] << 75) +
      (src075[42] << 75) +
      (src075[43] << 75) +
      (src075[44] << 75) +
      (src075[45] << 75) +
      (src075[46] << 75) +
      (src075[47] << 75) +
      (src075[48] << 75) +
      (src075[49] << 75) +
      (src075[50] << 75) +
      (src075[51] << 75) +
      (src076[0] << 76) +
      (src076[1] << 76) +
      (src076[2] << 76) +
      (src076[3] << 76) +
      (src076[4] << 76) +
      (src076[5] << 76) +
      (src076[6] << 76) +
      (src076[7] << 76) +
      (src076[8] << 76) +
      (src076[9] << 76) +
      (src076[10] << 76) +
      (src076[11] << 76) +
      (src076[12] << 76) +
      (src076[13] << 76) +
      (src076[14] << 76) +
      (src076[15] << 76) +
      (src076[16] << 76) +
      (src076[17] << 76) +
      (src076[18] << 76) +
      (src076[19] << 76) +
      (src076[20] << 76) +
      (src076[21] << 76) +
      (src076[22] << 76) +
      (src076[23] << 76) +
      (src076[24] << 76) +
      (src076[25] << 76) +
      (src076[26] << 76) +
      (src076[27] << 76) +
      (src076[28] << 76) +
      (src076[29] << 76) +
      (src076[30] << 76) +
      (src076[31] << 76) +
      (src076[32] << 76) +
      (src076[33] << 76) +
      (src076[34] << 76) +
      (src076[35] << 76) +
      (src076[36] << 76) +
      (src076[37] << 76) +
      (src076[38] << 76) +
      (src076[39] << 76) +
      (src076[40] << 76) +
      (src076[41] << 76) +
      (src076[42] << 76) +
      (src076[43] << 76) +
      (src076[44] << 76) +
      (src076[45] << 76) +
      (src076[46] << 76) +
      (src076[47] << 76) +
      (src076[48] << 76) +
      (src076[49] << 76) +
      (src076[50] << 76) +
      (src077[0] << 77) +
      (src077[1] << 77) +
      (src077[2] << 77) +
      (src077[3] << 77) +
      (src077[4] << 77) +
      (src077[5] << 77) +
      (src077[6] << 77) +
      (src077[7] << 77) +
      (src077[8] << 77) +
      (src077[9] << 77) +
      (src077[10] << 77) +
      (src077[11] << 77) +
      (src077[12] << 77) +
      (src077[13] << 77) +
      (src077[14] << 77) +
      (src077[15] << 77) +
      (src077[16] << 77) +
      (src077[17] << 77) +
      (src077[18] << 77) +
      (src077[19] << 77) +
      (src077[20] << 77) +
      (src077[21] << 77) +
      (src077[22] << 77) +
      (src077[23] << 77) +
      (src077[24] << 77) +
      (src077[25] << 77) +
      (src077[26] << 77) +
      (src077[27] << 77) +
      (src077[28] << 77) +
      (src077[29] << 77) +
      (src077[30] << 77) +
      (src077[31] << 77) +
      (src077[32] << 77) +
      (src077[33] << 77) +
      (src077[34] << 77) +
      (src077[35] << 77) +
      (src077[36] << 77) +
      (src077[37] << 77) +
      (src077[38] << 77) +
      (src077[39] << 77) +
      (src077[40] << 77) +
      (src077[41] << 77) +
      (src077[42] << 77) +
      (src077[43] << 77) +
      (src077[44] << 77) +
      (src077[45] << 77) +
      (src077[46] << 77) +
      (src077[47] << 77) +
      (src077[48] << 77) +
      (src077[49] << 77) +
      (src078[0] << 78) +
      (src078[1] << 78) +
      (src078[2] << 78) +
      (src078[3] << 78) +
      (src078[4] << 78) +
      (src078[5] << 78) +
      (src078[6] << 78) +
      (src078[7] << 78) +
      (src078[8] << 78) +
      (src078[9] << 78) +
      (src078[10] << 78) +
      (src078[11] << 78) +
      (src078[12] << 78) +
      (src078[13] << 78) +
      (src078[14] << 78) +
      (src078[15] << 78) +
      (src078[16] << 78) +
      (src078[17] << 78) +
      (src078[18] << 78) +
      (src078[19] << 78) +
      (src078[20] << 78) +
      (src078[21] << 78) +
      (src078[22] << 78) +
      (src078[23] << 78) +
      (src078[24] << 78) +
      (src078[25] << 78) +
      (src078[26] << 78) +
      (src078[27] << 78) +
      (src078[28] << 78) +
      (src078[29] << 78) +
      (src078[30] << 78) +
      (src078[31] << 78) +
      (src078[32] << 78) +
      (src078[33] << 78) +
      (src078[34] << 78) +
      (src078[35] << 78) +
      (src078[36] << 78) +
      (src078[37] << 78) +
      (src078[38] << 78) +
      (src078[39] << 78) +
      (src078[40] << 78) +
      (src078[41] << 78) +
      (src078[42] << 78) +
      (src078[43] << 78) +
      (src078[44] << 78) +
      (src078[45] << 78) +
      (src078[46] << 78) +
      (src078[47] << 78) +
      (src078[48] << 78) +
      (src079[0] << 79) +
      (src079[1] << 79) +
      (src079[2] << 79) +
      (src079[3] << 79) +
      (src079[4] << 79) +
      (src079[5] << 79) +
      (src079[6] << 79) +
      (src079[7] << 79) +
      (src079[8] << 79) +
      (src079[9] << 79) +
      (src079[10] << 79) +
      (src079[11] << 79) +
      (src079[12] << 79) +
      (src079[13] << 79) +
      (src079[14] << 79) +
      (src079[15] << 79) +
      (src079[16] << 79) +
      (src079[17] << 79) +
      (src079[18] << 79) +
      (src079[19] << 79) +
      (src079[20] << 79) +
      (src079[21] << 79) +
      (src079[22] << 79) +
      (src079[23] << 79) +
      (src079[24] << 79) +
      (src079[25] << 79) +
      (src079[26] << 79) +
      (src079[27] << 79) +
      (src079[28] << 79) +
      (src079[29] << 79) +
      (src079[30] << 79) +
      (src079[31] << 79) +
      (src079[32] << 79) +
      (src079[33] << 79) +
      (src079[34] << 79) +
      (src079[35] << 79) +
      (src079[36] << 79) +
      (src079[37] << 79) +
      (src079[38] << 79) +
      (src079[39] << 79) +
      (src079[40] << 79) +
      (src079[41] << 79) +
      (src079[42] << 79) +
      (src079[43] << 79) +
      (src079[44] << 79) +
      (src079[45] << 79) +
      (src079[46] << 79) +
      (src079[47] << 79) +
      (src080[0] << 80) +
      (src080[1] << 80) +
      (src080[2] << 80) +
      (src080[3] << 80) +
      (src080[4] << 80) +
      (src080[5] << 80) +
      (src080[6] << 80) +
      (src080[7] << 80) +
      (src080[8] << 80) +
      (src080[9] << 80) +
      (src080[10] << 80) +
      (src080[11] << 80) +
      (src080[12] << 80) +
      (src080[13] << 80) +
      (src080[14] << 80) +
      (src080[15] << 80) +
      (src080[16] << 80) +
      (src080[17] << 80) +
      (src080[18] << 80) +
      (src080[19] << 80) +
      (src080[20] << 80) +
      (src080[21] << 80) +
      (src080[22] << 80) +
      (src080[23] << 80) +
      (src080[24] << 80) +
      (src080[25] << 80) +
      (src080[26] << 80) +
      (src080[27] << 80) +
      (src080[28] << 80) +
      (src080[29] << 80) +
      (src080[30] << 80) +
      (src080[31] << 80) +
      (src080[32] << 80) +
      (src080[33] << 80) +
      (src080[34] << 80) +
      (src080[35] << 80) +
      (src080[36] << 80) +
      (src080[37] << 80) +
      (src080[38] << 80) +
      (src080[39] << 80) +
      (src080[40] << 80) +
      (src080[41] << 80) +
      (src080[42] << 80) +
      (src080[43] << 80) +
      (src080[44] << 80) +
      (src080[45] << 80) +
      (src080[46] << 80) +
      (src081[0] << 81) +
      (src081[1] << 81) +
      (src081[2] << 81) +
      (src081[3] << 81) +
      (src081[4] << 81) +
      (src081[5] << 81) +
      (src081[6] << 81) +
      (src081[7] << 81) +
      (src081[8] << 81) +
      (src081[9] << 81) +
      (src081[10] << 81) +
      (src081[11] << 81) +
      (src081[12] << 81) +
      (src081[13] << 81) +
      (src081[14] << 81) +
      (src081[15] << 81) +
      (src081[16] << 81) +
      (src081[17] << 81) +
      (src081[18] << 81) +
      (src081[19] << 81) +
      (src081[20] << 81) +
      (src081[21] << 81) +
      (src081[22] << 81) +
      (src081[23] << 81) +
      (src081[24] << 81) +
      (src081[25] << 81) +
      (src081[26] << 81) +
      (src081[27] << 81) +
      (src081[28] << 81) +
      (src081[29] << 81) +
      (src081[30] << 81) +
      (src081[31] << 81) +
      (src081[32] << 81) +
      (src081[33] << 81) +
      (src081[34] << 81) +
      (src081[35] << 81) +
      (src081[36] << 81) +
      (src081[37] << 81) +
      (src081[38] << 81) +
      (src081[39] << 81) +
      (src081[40] << 81) +
      (src081[41] << 81) +
      (src081[42] << 81) +
      (src081[43] << 81) +
      (src081[44] << 81) +
      (src081[45] << 81) +
      (src082[0] << 82) +
      (src082[1] << 82) +
      (src082[2] << 82) +
      (src082[3] << 82) +
      (src082[4] << 82) +
      (src082[5] << 82) +
      (src082[6] << 82) +
      (src082[7] << 82) +
      (src082[8] << 82) +
      (src082[9] << 82) +
      (src082[10] << 82) +
      (src082[11] << 82) +
      (src082[12] << 82) +
      (src082[13] << 82) +
      (src082[14] << 82) +
      (src082[15] << 82) +
      (src082[16] << 82) +
      (src082[17] << 82) +
      (src082[18] << 82) +
      (src082[19] << 82) +
      (src082[20] << 82) +
      (src082[21] << 82) +
      (src082[22] << 82) +
      (src082[23] << 82) +
      (src082[24] << 82) +
      (src082[25] << 82) +
      (src082[26] << 82) +
      (src082[27] << 82) +
      (src082[28] << 82) +
      (src082[29] << 82) +
      (src082[30] << 82) +
      (src082[31] << 82) +
      (src082[32] << 82) +
      (src082[33] << 82) +
      (src082[34] << 82) +
      (src082[35] << 82) +
      (src082[36] << 82) +
      (src082[37] << 82) +
      (src082[38] << 82) +
      (src082[39] << 82) +
      (src082[40] << 82) +
      (src082[41] << 82) +
      (src082[42] << 82) +
      (src082[43] << 82) +
      (src082[44] << 82) +
      (src083[0] << 83) +
      (src083[1] << 83) +
      (src083[2] << 83) +
      (src083[3] << 83) +
      (src083[4] << 83) +
      (src083[5] << 83) +
      (src083[6] << 83) +
      (src083[7] << 83) +
      (src083[8] << 83) +
      (src083[9] << 83) +
      (src083[10] << 83) +
      (src083[11] << 83) +
      (src083[12] << 83) +
      (src083[13] << 83) +
      (src083[14] << 83) +
      (src083[15] << 83) +
      (src083[16] << 83) +
      (src083[17] << 83) +
      (src083[18] << 83) +
      (src083[19] << 83) +
      (src083[20] << 83) +
      (src083[21] << 83) +
      (src083[22] << 83) +
      (src083[23] << 83) +
      (src083[24] << 83) +
      (src083[25] << 83) +
      (src083[26] << 83) +
      (src083[27] << 83) +
      (src083[28] << 83) +
      (src083[29] << 83) +
      (src083[30] << 83) +
      (src083[31] << 83) +
      (src083[32] << 83) +
      (src083[33] << 83) +
      (src083[34] << 83) +
      (src083[35] << 83) +
      (src083[36] << 83) +
      (src083[37] << 83) +
      (src083[38] << 83) +
      (src083[39] << 83) +
      (src083[40] << 83) +
      (src083[41] << 83) +
      (src083[42] << 83) +
      (src083[43] << 83) +
      (src084[0] << 84) +
      (src084[1] << 84) +
      (src084[2] << 84) +
      (src084[3] << 84) +
      (src084[4] << 84) +
      (src084[5] << 84) +
      (src084[6] << 84) +
      (src084[7] << 84) +
      (src084[8] << 84) +
      (src084[9] << 84) +
      (src084[10] << 84) +
      (src084[11] << 84) +
      (src084[12] << 84) +
      (src084[13] << 84) +
      (src084[14] << 84) +
      (src084[15] << 84) +
      (src084[16] << 84) +
      (src084[17] << 84) +
      (src084[18] << 84) +
      (src084[19] << 84) +
      (src084[20] << 84) +
      (src084[21] << 84) +
      (src084[22] << 84) +
      (src084[23] << 84) +
      (src084[24] << 84) +
      (src084[25] << 84) +
      (src084[26] << 84) +
      (src084[27] << 84) +
      (src084[28] << 84) +
      (src084[29] << 84) +
      (src084[30] << 84) +
      (src084[31] << 84) +
      (src084[32] << 84) +
      (src084[33] << 84) +
      (src084[34] << 84) +
      (src084[35] << 84) +
      (src084[36] << 84) +
      (src084[37] << 84) +
      (src084[38] << 84) +
      (src084[39] << 84) +
      (src084[40] << 84) +
      (src084[41] << 84) +
      (src084[42] << 84) +
      (src085[0] << 85) +
      (src085[1] << 85) +
      (src085[2] << 85) +
      (src085[3] << 85) +
      (src085[4] << 85) +
      (src085[5] << 85) +
      (src085[6] << 85) +
      (src085[7] << 85) +
      (src085[8] << 85) +
      (src085[9] << 85) +
      (src085[10] << 85) +
      (src085[11] << 85) +
      (src085[12] << 85) +
      (src085[13] << 85) +
      (src085[14] << 85) +
      (src085[15] << 85) +
      (src085[16] << 85) +
      (src085[17] << 85) +
      (src085[18] << 85) +
      (src085[19] << 85) +
      (src085[20] << 85) +
      (src085[21] << 85) +
      (src085[22] << 85) +
      (src085[23] << 85) +
      (src085[24] << 85) +
      (src085[25] << 85) +
      (src085[26] << 85) +
      (src085[27] << 85) +
      (src085[28] << 85) +
      (src085[29] << 85) +
      (src085[30] << 85) +
      (src085[31] << 85) +
      (src085[32] << 85) +
      (src085[33] << 85) +
      (src085[34] << 85) +
      (src085[35] << 85) +
      (src085[36] << 85) +
      (src085[37] << 85) +
      (src085[38] << 85) +
      (src085[39] << 85) +
      (src085[40] << 85) +
      (src085[41] << 85) +
      (src086[0] << 86) +
      (src086[1] << 86) +
      (src086[2] << 86) +
      (src086[3] << 86) +
      (src086[4] << 86) +
      (src086[5] << 86) +
      (src086[6] << 86) +
      (src086[7] << 86) +
      (src086[8] << 86) +
      (src086[9] << 86) +
      (src086[10] << 86) +
      (src086[11] << 86) +
      (src086[12] << 86) +
      (src086[13] << 86) +
      (src086[14] << 86) +
      (src086[15] << 86) +
      (src086[16] << 86) +
      (src086[17] << 86) +
      (src086[18] << 86) +
      (src086[19] << 86) +
      (src086[20] << 86) +
      (src086[21] << 86) +
      (src086[22] << 86) +
      (src086[23] << 86) +
      (src086[24] << 86) +
      (src086[25] << 86) +
      (src086[26] << 86) +
      (src086[27] << 86) +
      (src086[28] << 86) +
      (src086[29] << 86) +
      (src086[30] << 86) +
      (src086[31] << 86) +
      (src086[32] << 86) +
      (src086[33] << 86) +
      (src086[34] << 86) +
      (src086[35] << 86) +
      (src086[36] << 86) +
      (src086[37] << 86) +
      (src086[38] << 86) +
      (src086[39] << 86) +
      (src086[40] << 86) +
      (src087[0] << 87) +
      (src087[1] << 87) +
      (src087[2] << 87) +
      (src087[3] << 87) +
      (src087[4] << 87) +
      (src087[5] << 87) +
      (src087[6] << 87) +
      (src087[7] << 87) +
      (src087[8] << 87) +
      (src087[9] << 87) +
      (src087[10] << 87) +
      (src087[11] << 87) +
      (src087[12] << 87) +
      (src087[13] << 87) +
      (src087[14] << 87) +
      (src087[15] << 87) +
      (src087[16] << 87) +
      (src087[17] << 87) +
      (src087[18] << 87) +
      (src087[19] << 87) +
      (src087[20] << 87) +
      (src087[21] << 87) +
      (src087[22] << 87) +
      (src087[23] << 87) +
      (src087[24] << 87) +
      (src087[25] << 87) +
      (src087[26] << 87) +
      (src087[27] << 87) +
      (src087[28] << 87) +
      (src087[29] << 87) +
      (src087[30] << 87) +
      (src087[31] << 87) +
      (src087[32] << 87) +
      (src087[33] << 87) +
      (src087[34] << 87) +
      (src087[35] << 87) +
      (src087[36] << 87) +
      (src087[37] << 87) +
      (src087[38] << 87) +
      (src087[39] << 87) +
      (src088[0] << 88) +
      (src088[1] << 88) +
      (src088[2] << 88) +
      (src088[3] << 88) +
      (src088[4] << 88) +
      (src088[5] << 88) +
      (src088[6] << 88) +
      (src088[7] << 88) +
      (src088[8] << 88) +
      (src088[9] << 88) +
      (src088[10] << 88) +
      (src088[11] << 88) +
      (src088[12] << 88) +
      (src088[13] << 88) +
      (src088[14] << 88) +
      (src088[15] << 88) +
      (src088[16] << 88) +
      (src088[17] << 88) +
      (src088[18] << 88) +
      (src088[19] << 88) +
      (src088[20] << 88) +
      (src088[21] << 88) +
      (src088[22] << 88) +
      (src088[23] << 88) +
      (src088[24] << 88) +
      (src088[25] << 88) +
      (src088[26] << 88) +
      (src088[27] << 88) +
      (src088[28] << 88) +
      (src088[29] << 88) +
      (src088[30] << 88) +
      (src088[31] << 88) +
      (src088[32] << 88) +
      (src088[33] << 88) +
      (src088[34] << 88) +
      (src088[35] << 88) +
      (src088[36] << 88) +
      (src088[37] << 88) +
      (src088[38] << 88) +
      (src089[0] << 89) +
      (src089[1] << 89) +
      (src089[2] << 89) +
      (src089[3] << 89) +
      (src089[4] << 89) +
      (src089[5] << 89) +
      (src089[6] << 89) +
      (src089[7] << 89) +
      (src089[8] << 89) +
      (src089[9] << 89) +
      (src089[10] << 89) +
      (src089[11] << 89) +
      (src089[12] << 89) +
      (src089[13] << 89) +
      (src089[14] << 89) +
      (src089[15] << 89) +
      (src089[16] << 89) +
      (src089[17] << 89) +
      (src089[18] << 89) +
      (src089[19] << 89) +
      (src089[20] << 89) +
      (src089[21] << 89) +
      (src089[22] << 89) +
      (src089[23] << 89) +
      (src089[24] << 89) +
      (src089[25] << 89) +
      (src089[26] << 89) +
      (src089[27] << 89) +
      (src089[28] << 89) +
      (src089[29] << 89) +
      (src089[30] << 89) +
      (src089[31] << 89) +
      (src089[32] << 89) +
      (src089[33] << 89) +
      (src089[34] << 89) +
      (src089[35] << 89) +
      (src089[36] << 89) +
      (src089[37] << 89) +
      (src090[0] << 90) +
      (src090[1] << 90) +
      (src090[2] << 90) +
      (src090[3] << 90) +
      (src090[4] << 90) +
      (src090[5] << 90) +
      (src090[6] << 90) +
      (src090[7] << 90) +
      (src090[8] << 90) +
      (src090[9] << 90) +
      (src090[10] << 90) +
      (src090[11] << 90) +
      (src090[12] << 90) +
      (src090[13] << 90) +
      (src090[14] << 90) +
      (src090[15] << 90) +
      (src090[16] << 90) +
      (src090[17] << 90) +
      (src090[18] << 90) +
      (src090[19] << 90) +
      (src090[20] << 90) +
      (src090[21] << 90) +
      (src090[22] << 90) +
      (src090[23] << 90) +
      (src090[24] << 90) +
      (src090[25] << 90) +
      (src090[26] << 90) +
      (src090[27] << 90) +
      (src090[28] << 90) +
      (src090[29] << 90) +
      (src090[30] << 90) +
      (src090[31] << 90) +
      (src090[32] << 90) +
      (src090[33] << 90) +
      (src090[34] << 90) +
      (src090[35] << 90) +
      (src090[36] << 90) +
      (src091[0] << 91) +
      (src091[1] << 91) +
      (src091[2] << 91) +
      (src091[3] << 91) +
      (src091[4] << 91) +
      (src091[5] << 91) +
      (src091[6] << 91) +
      (src091[7] << 91) +
      (src091[8] << 91) +
      (src091[9] << 91) +
      (src091[10] << 91) +
      (src091[11] << 91) +
      (src091[12] << 91) +
      (src091[13] << 91) +
      (src091[14] << 91) +
      (src091[15] << 91) +
      (src091[16] << 91) +
      (src091[17] << 91) +
      (src091[18] << 91) +
      (src091[19] << 91) +
      (src091[20] << 91) +
      (src091[21] << 91) +
      (src091[22] << 91) +
      (src091[23] << 91) +
      (src091[24] << 91) +
      (src091[25] << 91) +
      (src091[26] << 91) +
      (src091[27] << 91) +
      (src091[28] << 91) +
      (src091[29] << 91) +
      (src091[30] << 91) +
      (src091[31] << 91) +
      (src091[32] << 91) +
      (src091[33] << 91) +
      (src091[34] << 91) +
      (src091[35] << 91) +
      (src092[0] << 92) +
      (src092[1] << 92) +
      (src092[2] << 92) +
      (src092[3] << 92) +
      (src092[4] << 92) +
      (src092[5] << 92) +
      (src092[6] << 92) +
      (src092[7] << 92) +
      (src092[8] << 92) +
      (src092[9] << 92) +
      (src092[10] << 92) +
      (src092[11] << 92) +
      (src092[12] << 92) +
      (src092[13] << 92) +
      (src092[14] << 92) +
      (src092[15] << 92) +
      (src092[16] << 92) +
      (src092[17] << 92) +
      (src092[18] << 92) +
      (src092[19] << 92) +
      (src092[20] << 92) +
      (src092[21] << 92) +
      (src092[22] << 92) +
      (src092[23] << 92) +
      (src092[24] << 92) +
      (src092[25] << 92) +
      (src092[26] << 92) +
      (src092[27] << 92) +
      (src092[28] << 92) +
      (src092[29] << 92) +
      (src092[30] << 92) +
      (src092[31] << 92) +
      (src092[32] << 92) +
      (src092[33] << 92) +
      (src092[34] << 92) +
      (src093[0] << 93) +
      (src093[1] << 93) +
      (src093[2] << 93) +
      (src093[3] << 93) +
      (src093[4] << 93) +
      (src093[5] << 93) +
      (src093[6] << 93) +
      (src093[7] << 93) +
      (src093[8] << 93) +
      (src093[9] << 93) +
      (src093[10] << 93) +
      (src093[11] << 93) +
      (src093[12] << 93) +
      (src093[13] << 93) +
      (src093[14] << 93) +
      (src093[15] << 93) +
      (src093[16] << 93) +
      (src093[17] << 93) +
      (src093[18] << 93) +
      (src093[19] << 93) +
      (src093[20] << 93) +
      (src093[21] << 93) +
      (src093[22] << 93) +
      (src093[23] << 93) +
      (src093[24] << 93) +
      (src093[25] << 93) +
      (src093[26] << 93) +
      (src093[27] << 93) +
      (src093[28] << 93) +
      (src093[29] << 93) +
      (src093[30] << 93) +
      (src093[31] << 93) +
      (src093[32] << 93) +
      (src093[33] << 93) +
      (src094[0] << 94) +
      (src094[1] << 94) +
      (src094[2] << 94) +
      (src094[3] << 94) +
      (src094[4] << 94) +
      (src094[5] << 94) +
      (src094[6] << 94) +
      (src094[7] << 94) +
      (src094[8] << 94) +
      (src094[9] << 94) +
      (src094[10] << 94) +
      (src094[11] << 94) +
      (src094[12] << 94) +
      (src094[13] << 94) +
      (src094[14] << 94) +
      (src094[15] << 94) +
      (src094[16] << 94) +
      (src094[17] << 94) +
      (src094[18] << 94) +
      (src094[19] << 94) +
      (src094[20] << 94) +
      (src094[21] << 94) +
      (src094[22] << 94) +
      (src094[23] << 94) +
      (src094[24] << 94) +
      (src094[25] << 94) +
      (src094[26] << 94) +
      (src094[27] << 94) +
      (src094[28] << 94) +
      (src094[29] << 94) +
      (src094[30] << 94) +
      (src094[31] << 94) +
      (src094[32] << 94) +
      (src095[0] << 95) +
      (src095[1] << 95) +
      (src095[2] << 95) +
      (src095[3] << 95) +
      (src095[4] << 95) +
      (src095[5] << 95) +
      (src095[6] << 95) +
      (src095[7] << 95) +
      (src095[8] << 95) +
      (src095[9] << 95) +
      (src095[10] << 95) +
      (src095[11] << 95) +
      (src095[12] << 95) +
      (src095[13] << 95) +
      (src095[14] << 95) +
      (src095[15] << 95) +
      (src095[16] << 95) +
      (src095[17] << 95) +
      (src095[18] << 95) +
      (src095[19] << 95) +
      (src095[20] << 95) +
      (src095[21] << 95) +
      (src095[22] << 95) +
      (src095[23] << 95) +
      (src095[24] << 95) +
      (src095[25] << 95) +
      (src095[26] << 95) +
      (src095[27] << 95) +
      (src095[28] << 95) +
      (src095[29] << 95) +
      (src095[30] << 95) +
      (src095[31] << 95) +
      (src096[0] << 96) +
      (src096[1] << 96) +
      (src096[2] << 96) +
      (src096[3] << 96) +
      (src096[4] << 96) +
      (src096[5] << 96) +
      (src096[6] << 96) +
      (src096[7] << 96) +
      (src096[8] << 96) +
      (src096[9] << 96) +
      (src096[10] << 96) +
      (src096[11] << 96) +
      (src096[12] << 96) +
      (src096[13] << 96) +
      (src096[14] << 96) +
      (src096[15] << 96) +
      (src096[16] << 96) +
      (src096[17] << 96) +
      (src096[18] << 96) +
      (src096[19] << 96) +
      (src096[20] << 96) +
      (src096[21] << 96) +
      (src096[22] << 96) +
      (src096[23] << 96) +
      (src096[24] << 96) +
      (src096[25] << 96) +
      (src096[26] << 96) +
      (src096[27] << 96) +
      (src096[28] << 96) +
      (src096[29] << 96) +
      (src096[30] << 96) +
      (src097[0] << 97) +
      (src097[1] << 97) +
      (src097[2] << 97) +
      (src097[3] << 97) +
      (src097[4] << 97) +
      (src097[5] << 97) +
      (src097[6] << 97) +
      (src097[7] << 97) +
      (src097[8] << 97) +
      (src097[9] << 97) +
      (src097[10] << 97) +
      (src097[11] << 97) +
      (src097[12] << 97) +
      (src097[13] << 97) +
      (src097[14] << 97) +
      (src097[15] << 97) +
      (src097[16] << 97) +
      (src097[17] << 97) +
      (src097[18] << 97) +
      (src097[19] << 97) +
      (src097[20] << 97) +
      (src097[21] << 97) +
      (src097[22] << 97) +
      (src097[23] << 97) +
      (src097[24] << 97) +
      (src097[25] << 97) +
      (src097[26] << 97) +
      (src097[27] << 97) +
      (src097[28] << 97) +
      (src097[29] << 97) +
      (src098[0] << 98) +
      (src098[1] << 98) +
      (src098[2] << 98) +
      (src098[3] << 98) +
      (src098[4] << 98) +
      (src098[5] << 98) +
      (src098[6] << 98) +
      (src098[7] << 98) +
      (src098[8] << 98) +
      (src098[9] << 98) +
      (src098[10] << 98) +
      (src098[11] << 98) +
      (src098[12] << 98) +
      (src098[13] << 98) +
      (src098[14] << 98) +
      (src098[15] << 98) +
      (src098[16] << 98) +
      (src098[17] << 98) +
      (src098[18] << 98) +
      (src098[19] << 98) +
      (src098[20] << 98) +
      (src098[21] << 98) +
      (src098[22] << 98) +
      (src098[23] << 98) +
      (src098[24] << 98) +
      (src098[25] << 98) +
      (src098[26] << 98) +
      (src098[27] << 98) +
      (src098[28] << 98) +
      (src099[0] << 99) +
      (src099[1] << 99) +
      (src099[2] << 99) +
      (src099[3] << 99) +
      (src099[4] << 99) +
      (src099[5] << 99) +
      (src099[6] << 99) +
      (src099[7] << 99) +
      (src099[8] << 99) +
      (src099[9] << 99) +
      (src099[10] << 99) +
      (src099[11] << 99) +
      (src099[12] << 99) +
      (src099[13] << 99) +
      (src099[14] << 99) +
      (src099[15] << 99) +
      (src099[16] << 99) +
      (src099[17] << 99) +
      (src099[18] << 99) +
      (src099[19] << 99) +
      (src099[20] << 99) +
      (src099[21] << 99) +
      (src099[22] << 99) +
      (src099[23] << 99) +
      (src099[24] << 99) +
      (src099[25] << 99) +
      (src099[26] << 99) +
      (src099[27] << 99) +
      (src100[0] << 100) +
      (src100[1] << 100) +
      (src100[2] << 100) +
      (src100[3] << 100) +
      (src100[4] << 100) +
      (src100[5] << 100) +
      (src100[6] << 100) +
      (src100[7] << 100) +
      (src100[8] << 100) +
      (src100[9] << 100) +
      (src100[10] << 100) +
      (src100[11] << 100) +
      (src100[12] << 100) +
      (src100[13] << 100) +
      (src100[14] << 100) +
      (src100[15] << 100) +
      (src100[16] << 100) +
      (src100[17] << 100) +
      (src100[18] << 100) +
      (src100[19] << 100) +
      (src100[20] << 100) +
      (src100[21] << 100) +
      (src100[22] << 100) +
      (src100[23] << 100) +
      (src100[24] << 100) +
      (src100[25] << 100) +
      (src100[26] << 100) +
      (src101[0] << 101) +
      (src101[1] << 101) +
      (src101[2] << 101) +
      (src101[3] << 101) +
      (src101[4] << 101) +
      (src101[5] << 101) +
      (src101[6] << 101) +
      (src101[7] << 101) +
      (src101[8] << 101) +
      (src101[9] << 101) +
      (src101[10] << 101) +
      (src101[11] << 101) +
      (src101[12] << 101) +
      (src101[13] << 101) +
      (src101[14] << 101) +
      (src101[15] << 101) +
      (src101[16] << 101) +
      (src101[17] << 101) +
      (src101[18] << 101) +
      (src101[19] << 101) +
      (src101[20] << 101) +
      (src101[21] << 101) +
      (src101[22] << 101) +
      (src101[23] << 101) +
      (src101[24] << 101) +
      (src101[25] << 101) +
      (src102[0] << 102) +
      (src102[1] << 102) +
      (src102[2] << 102) +
      (src102[3] << 102) +
      (src102[4] << 102) +
      (src102[5] << 102) +
      (src102[6] << 102) +
      (src102[7] << 102) +
      (src102[8] << 102) +
      (src102[9] << 102) +
      (src102[10] << 102) +
      (src102[11] << 102) +
      (src102[12] << 102) +
      (src102[13] << 102) +
      (src102[14] << 102) +
      (src102[15] << 102) +
      (src102[16] << 102) +
      (src102[17] << 102) +
      (src102[18] << 102) +
      (src102[19] << 102) +
      (src102[20] << 102) +
      (src102[21] << 102) +
      (src102[22] << 102) +
      (src102[23] << 102) +
      (src102[24] << 102) +
      (src103[0] << 103) +
      (src103[1] << 103) +
      (src103[2] << 103) +
      (src103[3] << 103) +
      (src103[4] << 103) +
      (src103[5] << 103) +
      (src103[6] << 103) +
      (src103[7] << 103) +
      (src103[8] << 103) +
      (src103[9] << 103) +
      (src103[10] << 103) +
      (src103[11] << 103) +
      (src103[12] << 103) +
      (src103[13] << 103) +
      (src103[14] << 103) +
      (src103[15] << 103) +
      (src103[16] << 103) +
      (src103[17] << 103) +
      (src103[18] << 103) +
      (src103[19] << 103) +
      (src103[20] << 103) +
      (src103[21] << 103) +
      (src103[22] << 103) +
      (src103[23] << 103) +
      (src104[0] << 104) +
      (src104[1] << 104) +
      (src104[2] << 104) +
      (src104[3] << 104) +
      (src104[4] << 104) +
      (src104[5] << 104) +
      (src104[6] << 104) +
      (src104[7] << 104) +
      (src104[8] << 104) +
      (src104[9] << 104) +
      (src104[10] << 104) +
      (src104[11] << 104) +
      (src104[12] << 104) +
      (src104[13] << 104) +
      (src104[14] << 104) +
      (src104[15] << 104) +
      (src104[16] << 104) +
      (src104[17] << 104) +
      (src104[18] << 104) +
      (src104[19] << 104) +
      (src104[20] << 104) +
      (src104[21] << 104) +
      (src104[22] << 104) +
      (src105[0] << 105) +
      (src105[1] << 105) +
      (src105[2] << 105) +
      (src105[3] << 105) +
      (src105[4] << 105) +
      (src105[5] << 105) +
      (src105[6] << 105) +
      (src105[7] << 105) +
      (src105[8] << 105) +
      (src105[9] << 105) +
      (src105[10] << 105) +
      (src105[11] << 105) +
      (src105[12] << 105) +
      (src105[13] << 105) +
      (src105[14] << 105) +
      (src105[15] << 105) +
      (src105[16] << 105) +
      (src105[17] << 105) +
      (src105[18] << 105) +
      (src105[19] << 105) +
      (src105[20] << 105) +
      (src105[21] << 105) +
      (src106[0] << 106) +
      (src106[1] << 106) +
      (src106[2] << 106) +
      (src106[3] << 106) +
      (src106[4] << 106) +
      (src106[5] << 106) +
      (src106[6] << 106) +
      (src106[7] << 106) +
      (src106[8] << 106) +
      (src106[9] << 106) +
      (src106[10] << 106) +
      (src106[11] << 106) +
      (src106[12] << 106) +
      (src106[13] << 106) +
      (src106[14] << 106) +
      (src106[15] << 106) +
      (src106[16] << 106) +
      (src106[17] << 106) +
      (src106[18] << 106) +
      (src106[19] << 106) +
      (src106[20] << 106) +
      (src107[0] << 107) +
      (src107[1] << 107) +
      (src107[2] << 107) +
      (src107[3] << 107) +
      (src107[4] << 107) +
      (src107[5] << 107) +
      (src107[6] << 107) +
      (src107[7] << 107) +
      (src107[8] << 107) +
      (src107[9] << 107) +
      (src107[10] << 107) +
      (src107[11] << 107) +
      (src107[12] << 107) +
      (src107[13] << 107) +
      (src107[14] << 107) +
      (src107[15] << 107) +
      (src107[16] << 107) +
      (src107[17] << 107) +
      (src107[18] << 107) +
      (src107[19] << 107) +
      (src108[0] << 108) +
      (src108[1] << 108) +
      (src108[2] << 108) +
      (src108[3] << 108) +
      (src108[4] << 108) +
      (src108[5] << 108) +
      (src108[6] << 108) +
      (src108[7] << 108) +
      (src108[8] << 108) +
      (src108[9] << 108) +
      (src108[10] << 108) +
      (src108[11] << 108) +
      (src108[12] << 108) +
      (src108[13] << 108) +
      (src108[14] << 108) +
      (src108[15] << 108) +
      (src108[16] << 108) +
      (src108[17] << 108) +
      (src108[18] << 108) +
      (src109[0] << 109) +
      (src109[1] << 109) +
      (src109[2] << 109) +
      (src109[3] << 109) +
      (src109[4] << 109) +
      (src109[5] << 109) +
      (src109[6] << 109) +
      (src109[7] << 109) +
      (src109[8] << 109) +
      (src109[9] << 109) +
      (src109[10] << 109) +
      (src109[11] << 109) +
      (src109[12] << 109) +
      (src109[13] << 109) +
      (src109[14] << 109) +
      (src109[15] << 109) +
      (src109[16] << 109) +
      (src109[17] << 109) +
      (src110[0] << 110) +
      (src110[1] << 110) +
      (src110[2] << 110) +
      (src110[3] << 110) +
      (src110[4] << 110) +
      (src110[5] << 110) +
      (src110[6] << 110) +
      (src110[7] << 110) +
      (src110[8] << 110) +
      (src110[9] << 110) +
      (src110[10] << 110) +
      (src110[11] << 110) +
      (src110[12] << 110) +
      (src110[13] << 110) +
      (src110[14] << 110) +
      (src110[15] << 110) +
      (src110[16] << 110) +
      (src111[0] << 111) +
      (src111[1] << 111) +
      (src111[2] << 111) +
      (src111[3] << 111) +
      (src111[4] << 111) +
      (src111[5] << 111) +
      (src111[6] << 111) +
      (src111[7] << 111) +
      (src111[8] << 111) +
      (src111[9] << 111) +
      (src111[10] << 111) +
      (src111[11] << 111) +
      (src111[12] << 111) +
      (src111[13] << 111) +
      (src111[14] << 111) +
      (src111[15] << 111) +
      (src112[0] << 112) +
      (src112[1] << 112) +
      (src112[2] << 112) +
      (src112[3] << 112) +
      (src112[4] << 112) +
      (src112[5] << 112) +
      (src112[6] << 112) +
      (src112[7] << 112) +
      (src112[8] << 112) +
      (src112[9] << 112) +
      (src112[10] << 112) +
      (src112[11] << 112) +
      (src112[12] << 112) +
      (src112[13] << 112) +
      (src112[14] << 112) +
      (src113[0] << 113) +
      (src113[1] << 113) +
      (src113[2] << 113) +
      (src113[3] << 113) +
      (src113[4] << 113) +
      (src113[5] << 113) +
      (src113[6] << 113) +
      (src113[7] << 113) +
      (src113[8] << 113) +
      (src113[9] << 113) +
      (src113[10] << 113) +
      (src113[11] << 113) +
      (src113[12] << 113) +
      (src113[13] << 113) +
      (src114[0] << 114) +
      (src114[1] << 114) +
      (src114[2] << 114) +
      (src114[3] << 114) +
      (src114[4] << 114) +
      (src114[5] << 114) +
      (src114[6] << 114) +
      (src114[7] << 114) +
      (src114[8] << 114) +
      (src114[9] << 114) +
      (src114[10] << 114) +
      (src114[11] << 114) +
      (src114[12] << 114) +
      (src115[0] << 115) +
      (src115[1] << 115) +
      (src115[2] << 115) +
      (src115[3] << 115) +
      (src115[4] << 115) +
      (src115[5] << 115) +
      (src115[6] << 115) +
      (src115[7] << 115) +
      (src115[8] << 115) +
      (src115[9] << 115) +
      (src115[10] << 115) +
      (src115[11] << 115) +
      (src116[0] << 116) +
      (src116[1] << 116) +
      (src116[2] << 116) +
      (src116[3] << 116) +
      (src116[4] << 116) +
      (src116[5] << 116) +
      (src116[6] << 116) +
      (src116[7] << 116) +
      (src116[8] << 116) +
      (src116[9] << 116) +
      (src116[10] << 116) +
      (src117[0] << 117) +
      (src117[1] << 117) +
      (src117[2] << 117) +
      (src117[3] << 117) +
      (src117[4] << 117) +
      (src117[5] << 117) +
      (src117[6] << 117) +
      (src117[7] << 117) +
      (src117[8] << 117) +
      (src117[9] << 117) +
      (src118[0] << 118) +
      (src118[1] << 118) +
      (src118[2] << 118) +
      (src118[3] << 118) +
      (src118[4] << 118) +
      (src118[5] << 118) +
      (src118[6] << 118) +
      (src118[7] << 118) +
      (src118[8] << 118) +
      (src119[0] << 119) +
      (src119[1] << 119) +
      (src119[2] << 119) +
      (src119[3] << 119) +
      (src119[4] << 119) +
      (src119[5] << 119) +
      (src119[6] << 119) +
      (src119[7] << 119) +
      (src120[0] << 120) +
      (src120[1] << 120) +
      (src120[2] << 120) +
      (src120[3] << 120) +
      (src120[4] << 120) +
      (src120[5] << 120) +
      (src120[6] << 120) +
      (src121[0] << 121) +
      (src121[1] << 121) +
      (src121[2] << 121) +
      (src121[3] << 121) +
      (src121[4] << 121) +
      (src121[5] << 121) +
      (src122[0] << 122) +
      (src122[1] << 122) +
      (src122[2] << 122) +
      (src122[3] << 122) +
      (src122[4] << 122) +
      (src123[0] << 123) +
      (src123[1] << 123) +
      (src123[2] << 123) +
      (src123[3] << 123) +
      (src124[0] << 124) +
      (src124[1] << 124) +
      (src124[2] << 124) +
      (src125[0] << 125) +
      (src125[1] << 125) +
      (src126[0] << 126);
   assign dstsum =
      (dst000[0] << 0) +
      (dst001[0] << 1) +
      (dst002[0] << 2) +
      (dst003[0] << 3) +
      (dst004[0] << 4) +
      (dst005[0] << 5) +
      (dst005[1] << 5) +
      (dst006[0] << 6) +
      (dst006[1] << 6) +
      (dst007[0] << 7) +
      (dst008[0] << 8) +
      (dst009[0] << 9) +
      (dst009[1] << 9) +
      (dst010[0] << 10) +
      (dst010[1] << 10) +
      (dst011[0] << 11) +
      (dst011[1] << 11) +
      (dst012[0] << 12) +
      (dst013[0] << 13) +
      (dst013[1] << 13) +
      (dst014[0] << 14) +
      (dst014[1] << 14) +
      (dst015[0] << 15) +
      (dst015[1] << 15) +
      (dst016[0] << 16) +
      (dst016[1] << 16) +
      (dst017[0] << 17) +
      (dst017[1] << 17) +
      (dst018[0] << 18) +
      (dst018[1] << 18) +
      (dst019[0] << 19) +
      (dst019[1] << 19) +
      (dst020[0] << 20) +
      (dst020[1] << 20) +
      (dst021[0] << 21) +
      (dst022[0] << 22) +
      (dst022[1] << 22) +
      (dst023[0] << 23) +
      (dst023[1] << 23) +
      (dst024[0] << 24) +
      (dst025[0] << 25) +
      (dst025[1] << 25) +
      (dst026[0] << 26) +
      (dst026[1] << 26) +
      (dst027[0] << 27) +
      (dst027[1] << 27) +
      (dst028[0] << 28) +
      (dst028[1] << 28) +
      (dst029[0] << 29) +
      (dst029[1] << 29) +
      (dst030[0] << 30) +
      (dst030[1] << 30) +
      (dst031[0] << 31) +
      (dst031[1] << 31) +
      (dst032[0] << 32) +
      (dst032[1] << 32) +
      (dst033[0] << 33) +
      (dst033[1] << 33) +
      (dst034[0] << 34) +
      (dst034[1] << 34) +
      (dst035[0] << 35) +
      (dst035[1] << 35) +
      (dst036[0] << 36) +
      (dst037[0] << 37) +
      (dst037[1] << 37) +
      (dst038[0] << 38) +
      (dst038[1] << 38) +
      (dst039[0] << 39) +
      (dst039[1] << 39) +
      (dst040[0] << 40) +
      (dst040[1] << 40) +
      (dst041[0] << 41) +
      (dst041[1] << 41) +
      (dst042[0] << 42) +
      (dst042[1] << 42) +
      (dst043[0] << 43) +
      (dst043[1] << 43) +
      (dst044[0] << 44) +
      (dst044[1] << 44) +
      (dst045[0] << 45) +
      (dst045[1] << 45) +
      (dst046[0] << 46) +
      (dst046[1] << 46) +
      (dst047[0] << 47) +
      (dst047[1] << 47) +
      (dst048[0] << 48) +
      (dst048[1] << 48) +
      (dst049[0] << 49) +
      (dst049[1] << 49) +
      (dst050[0] << 50) +
      (dst050[1] << 50) +
      (dst051[0] << 51) +
      (dst051[1] << 51) +
      (dst052[0] << 52) +
      (dst052[1] << 52) +
      (dst053[0] << 53) +
      (dst053[1] << 53) +
      (dst054[0] << 54) +
      (dst054[1] << 54) +
      (dst055[0] << 55) +
      (dst055[1] << 55) +
      (dst056[0] << 56) +
      (dst056[1] << 56) +
      (dst057[0] << 57) +
      (dst057[1] << 57) +
      (dst058[0] << 58) +
      (dst058[1] << 58) +
      (dst059[0] << 59) +
      (dst059[1] << 59) +
      (dst060[0] << 60) +
      (dst060[1] << 60) +
      (dst061[0] << 61) +
      (dst061[1] << 61) +
      (dst062[0] << 62) +
      (dst062[1] << 62) +
      (dst063[0] << 63) +
      (dst063[1] << 63) +
      (dst064[0] << 64) +
      (dst064[1] << 64) +
      (dst065[0] << 65) +
      (dst065[1] << 65) +
      (dst066[0] << 66) +
      (dst066[1] << 66) +
      (dst067[0] << 67) +
      (dst067[1] << 67) +
      (dst068[0] << 68) +
      (dst068[1] << 68) +
      (dst069[0] << 69) +
      (dst069[1] << 69) +
      (dst070[0] << 70) +
      (dst070[1] << 70) +
      (dst071[0] << 71) +
      (dst071[1] << 71) +
      (dst072[0] << 72) +
      (dst072[1] << 72) +
      (dst073[0] << 73) +
      (dst073[1] << 73) +
      (dst074[0] << 74) +
      (dst074[1] << 74) +
      (dst075[0] << 75) +
      (dst075[1] << 75) +
      (dst076[0] << 76) +
      (dst076[1] << 76) +
      (dst077[0] << 77) +
      (dst077[1] << 77) +
      (dst078[0] << 78) +
      (dst078[1] << 78) +
      (dst079[0] << 79) +
      (dst079[1] << 79) +
      (dst080[0] << 80) +
      (dst080[1] << 80) +
      (dst081[0] << 81) +
      (dst081[1] << 81) +
      (dst082[0] << 82) +
      (dst082[1] << 82) +
      (dst083[0] << 83) +
      (dst083[1] << 83) +
      (dst084[0] << 84) +
      (dst084[1] << 84) +
      (dst085[0] << 85) +
      (dst085[1] << 85) +
      (dst086[0] << 86) +
      (dst086[1] << 86) +
      (dst087[0] << 87) +
      (dst087[1] << 87) +
      (dst088[0] << 88) +
      (dst088[1] << 88) +
      (dst089[0] << 89) +
      (dst089[1] << 89) +
      (dst090[0] << 90) +
      (dst090[1] << 90) +
      (dst091[0] << 91) +
      (dst091[1] << 91) +
      (dst092[0] << 92) +
      (dst092[1] << 92) +
      (dst093[0] << 93) +
      (dst093[1] << 93) +
      (dst094[0] << 94) +
      (dst094[1] << 94) +
      (dst095[0] << 95) +
      (dst095[1] << 95) +
      (dst096[0] << 96) +
      (dst096[1] << 96) +
      (dst097[0] << 97) +
      (dst097[1] << 97) +
      (dst098[0] << 98) +
      (dst098[1] << 98) +
      (dst099[0] << 99) +
      (dst099[1] << 99) +
      (dst100[0] << 100) +
      (dst100[1] << 100) +
      (dst101[0] << 101) +
      (dst101[1] << 101) +
      (dst102[0] << 102) +
      (dst102[1] << 102) +
      (dst103[0] << 103) +
      (dst103[1] << 103) +
      (dst104[0] << 104) +
      (dst104[1] << 104) +
      (dst105[0] << 105) +
      (dst105[1] << 105) +
      (dst106[0] << 106) +
      (dst106[1] << 106) +
      (dst107[0] << 107) +
      (dst107[1] << 107) +
      (dst108[0] << 108) +
      (dst108[1] << 108) +
      (dst109[0] << 109) +
      (dst109[1] << 109) +
      (dst110[0] << 110) +
      (dst110[1] << 110) +
      (dst111[0] << 111) +
      (dst111[1] << 111) +
      (dst112[0] << 112) +
      (dst112[1] << 112) +
      (dst113[0] << 113) +
      (dst113[1] << 113) +
      (dst114[0] << 114) +
      (dst114[1] << 114) +
      (dst115[0] << 115) +
      (dst116[0] << 116) +
      (dst116[1] << 116) +
      (dst117[0] << 117) +
      (dst117[1] << 117) +
      (dst118[0] << 118) +
      (dst118[1] << 118) +
      (dst119[0] << 119) +
      (dst119[1] << 119) +
      (dst120[0] << 120) +
      (dst120[1] << 120) +
      (dst121[0] << 121) +
      (dst121[1] << 121) +
      (dst122[0] << 122) +
      (dst123[0] << 123) +
      (dst124[0] << 124) +
      (dst124[1] << 124) +
      (dst125[0] << 125) +
      (dst125[1] << 125) +
      (dst126[0] << 126) +
      (dst127[0] << 127) +
      (dst127[1] << 127) +
      (dst128[0] << 128);
   compressor main_cmp(src000, src001, src002, src003, src004, src005, src006, src007, src008, src009, src010, src011, src012, src013, src014, src015, src016, src017, src018, src019, src020, src021, src022, src023, src024, src025, src026, src027, src028, src029, src030, src031, src032, src033, src034, src035, src036, src037, src038, src039, src040, src041, src042, src043, src044, src045, src046, src047, src048, src049, src050, src051, src052, src053, src054, src055, src056, src057, src058, src059, src060, src061, src062, src063, src064, src065, src066, src067, src068, src069, src070, src071, src072, src073, src074, src075, src076, src077, src078, src079, src080, src081, src082, src083, src084, src085, src086, src087, src088, src089, src090, src091, src092, src093, src094, src095, src096, src097, src098, src099, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, dst000, dst001, dst002, dst003, dst004, dst005, dst006, dst007, dst008, dst009, dst010, dst011, dst012, dst013, dst014, dst015, dst016, dst017, dst018, dst019, dst020, dst021, dst022, dst023, dst024, dst025, dst026, dst027, dst028, dst029, dst030, dst031, dst032, dst033, dst034, dst035, dst036, dst037, dst038, dst039, dst040, dst041, dst042, dst043, dst044, dst045, dst046, dst047, dst048, dst049, dst050, dst051, dst052, dst053, dst054, dst055, dst056, dst057, dst058, dst059, dst060, dst061, dst062, dst063, dst064, dst065, dst066, dst067, dst068, dst069, dst070, dst071, dst072, dst073, dst074, dst075, dst076, dst077, dst078, dst079, dst080, dst081, dst082, dst083, dst084, dst085, dst086, dst087, dst088, dst089, dst090, dst091, dst092, dst093, dst094, dst095, dst096, dst097, dst098, dst099, dst100, dst101, dst102, dst103, dst104, dst105, dst106, dst107, dst108, dst109, dst110, dst111, dst112, dst113, dst114, dst115, dst116, dst117, dst118, dst119, dst120, dst121, dst122, dst123, dst124, dst125, dst126, dst127, dst128);
   assign test = srcsum == dstsum;
   initial begin
      $monitor("src: 0x%x, dst: 0x%x, test: %b", srcsum, dstsum, test);
   end
   initial begin
      src000 <= 1'h0;
      src001 <= 2'h0;
      src002 <= 3'h0;
      src003 <= 4'h0;
      src004 <= 5'h0;
      src005 <= 6'h0;
      src006 <= 7'h0;
      src007 <= 8'h0;
      src008 <= 9'h0;
      src009 <= 10'h0;
      src010 <= 11'h0;
      src011 <= 12'h0;
      src012 <= 13'h0;
      src013 <= 14'h0;
      src014 <= 15'h0;
      src015 <= 16'h0;
      src016 <= 17'h0;
      src017 <= 18'h0;
      src018 <= 19'h0;
      src019 <= 20'h0;
      src020 <= 21'h0;
      src021 <= 22'h0;
      src022 <= 23'h0;
      src023 <= 24'h0;
      src024 <= 25'h0;
      src025 <= 26'h0;
      src026 <= 27'h0;
      src027 <= 28'h0;
      src028 <= 29'h0;
      src029 <= 30'h0;
      src030 <= 31'h0;
      src031 <= 32'h0;
      src032 <= 33'h0;
      src033 <= 34'h0;
      src034 <= 35'h0;
      src035 <= 36'h0;
      src036 <= 37'h0;
      src037 <= 38'h0;
      src038 <= 39'h0;
      src039 <= 40'h0;
      src040 <= 41'h0;
      src041 <= 42'h0;
      src042 <= 43'h0;
      src043 <= 44'h0;
      src044 <= 45'h0;
      src045 <= 46'h0;
      src046 <= 47'h0;
      src047 <= 48'h0;
      src048 <= 49'h0;
      src049 <= 50'h0;
      src050 <= 51'h0;
      src051 <= 52'h0;
      src052 <= 53'h0;
      src053 <= 54'h0;
      src054 <= 55'h0;
      src055 <= 56'h0;
      src056 <= 57'h0;
      src057 <= 58'h0;
      src058 <= 59'h0;
      src059 <= 60'h0;
      src060 <= 61'h0;
      src061 <= 62'h0;
      src062 <= 63'h0;
      src063 <= 64'h0;
      src064 <= 63'h0;
      src065 <= 62'h0;
      src066 <= 61'h0;
      src067 <= 60'h0;
      src068 <= 59'h0;
      src069 <= 58'h0;
      src070 <= 57'h0;
      src071 <= 56'h0;
      src072 <= 55'h0;
      src073 <= 54'h0;
      src074 <= 53'h0;
      src075 <= 52'h0;
      src076 <= 51'h0;
      src077 <= 50'h0;
      src078 <= 49'h0;
      src079 <= 48'h0;
      src080 <= 47'h0;
      src081 <= 46'h0;
      src082 <= 45'h0;
      src083 <= 44'h0;
      src084 <= 43'h0;
      src085 <= 42'h0;
      src086 <= 41'h0;
      src087 <= 40'h0;
      src088 <= 39'h0;
      src089 <= 38'h0;
      src090 <= 37'h0;
      src091 <= 36'h0;
      src092 <= 35'h0;
      src093 <= 34'h0;
      src094 <= 33'h0;
      src095 <= 32'h0;
      src096 <= 31'h0;
      src097 <= 30'h0;
      src098 <= 29'h0;
      src099 <= 28'h0;
      src100 <= 27'h0;
      src101 <= 26'h0;
      src102 <= 25'h0;
      src103 <= 24'h0;
      src104 <= 23'h0;
      src105 <= 22'h0;
      src106 <= 21'h0;
      src107 <= 20'h0;
      src108 <= 19'h0;
      src109 <= 18'h0;
      src110 <= 17'h0;
      src111 <= 16'h0;
      src112 <= 15'h0;
      src113 <= 14'h0;
      src114 <= 13'h0;
      src115 <= 12'h0;
      src116 <= 11'h0;
      src117 <= 10'h0;
      src118 <= 9'h0;
      src119 <= 8'h0;
      src120 <= 7'h0;
      src121 <= 6'h0;
      src122 <= 5'h0;
      src123 <= 4'h0;
      src124 <= 3'h0;
      src125 <= 2'h0;
      src126 <= 1'h0;
      #1
      src000 <= 1'h1;
      src001 <= 2'h3;
      src002 <= 3'h7;
      src003 <= 4'hf;
      src004 <= 5'h1f;
      src005 <= 6'h3f;
      src006 <= 7'h7f;
      src007 <= 8'hff;
      src008 <= 9'h1ff;
      src009 <= 10'h3ff;
      src010 <= 11'h7ff;
      src011 <= 12'hfff;
      src012 <= 13'h1fff;
      src013 <= 14'h3fff;
      src014 <= 15'h7fff;
      src015 <= 16'hffff;
      src016 <= 17'h1ffff;
      src017 <= 18'h3ffff;
      src018 <= 19'h7ffff;
      src019 <= 20'hfffff;
      src020 <= 21'h1fffff;
      src021 <= 22'h3fffff;
      src022 <= 23'h7fffff;
      src023 <= 24'hffffff;
      src024 <= 25'h1ffffff;
      src025 <= 26'h3ffffff;
      src026 <= 27'h7ffffff;
      src027 <= 28'hfffffff;
      src028 <= 29'h1fffffff;
      src029 <= 30'h3fffffff;
      src030 <= 31'h7fffffff;
      src031 <= 32'hffffffff;
      src032 <= 33'h1ffffffff;
      src033 <= 34'h3ffffffff;
      src034 <= 35'h7ffffffff;
      src035 <= 36'hfffffffff;
      src036 <= 37'h1fffffffff;
      src037 <= 38'h3fffffffff;
      src038 <= 39'h7fffffffff;
      src039 <= 40'hffffffffff;
      src040 <= 41'h1ffffffffff;
      src041 <= 42'h3ffffffffff;
      src042 <= 43'h7ffffffffff;
      src043 <= 44'hfffffffffff;
      src044 <= 45'h1fffffffffff;
      src045 <= 46'h3fffffffffff;
      src046 <= 47'h7fffffffffff;
      src047 <= 48'hffffffffffff;
      src048 <= 49'h1ffffffffffff;
      src049 <= 50'h3ffffffffffff;
      src050 <= 51'h7ffffffffffff;
      src051 <= 52'hfffffffffffff;
      src052 <= 53'h1fffffffffffff;
      src053 <= 54'h3fffffffffffff;
      src054 <= 55'h7fffffffffffff;
      src055 <= 56'hffffffffffffff;
      src056 <= 57'h1ffffffffffffff;
      src057 <= 58'h3ffffffffffffff;
      src058 <= 59'h7ffffffffffffff;
      src059 <= 60'hfffffffffffffff;
      src060 <= 61'h1fffffffffffffff;
      src061 <= 62'h3fffffffffffffff;
      src062 <= 63'h7fffffffffffffff;
      src063 <= 64'hffffffffffffffff;
      src064 <= 63'h7fffffffffffffff;
      src065 <= 62'h3fffffffffffffff;
      src066 <= 61'h1fffffffffffffff;
      src067 <= 60'hfffffffffffffff;
      src068 <= 59'h7ffffffffffffff;
      src069 <= 58'h3ffffffffffffff;
      src070 <= 57'h1ffffffffffffff;
      src071 <= 56'hffffffffffffff;
      src072 <= 55'h7fffffffffffff;
      src073 <= 54'h3fffffffffffff;
      src074 <= 53'h1fffffffffffff;
      src075 <= 52'hfffffffffffff;
      src076 <= 51'h7ffffffffffff;
      src077 <= 50'h3ffffffffffff;
      src078 <= 49'h1ffffffffffff;
      src079 <= 48'hffffffffffff;
      src080 <= 47'h7fffffffffff;
      src081 <= 46'h3fffffffffff;
      src082 <= 45'h1fffffffffff;
      src083 <= 44'hfffffffffff;
      src084 <= 43'h7ffffffffff;
      src085 <= 42'h3ffffffffff;
      src086 <= 41'h1ffffffffff;
      src087 <= 40'hffffffffff;
      src088 <= 39'h7fffffffff;
      src089 <= 38'h3fffffffff;
      src090 <= 37'h1fffffffff;
      src091 <= 36'hfffffffff;
      src092 <= 35'h7ffffffff;
      src093 <= 34'h3ffffffff;
      src094 <= 33'h1ffffffff;
      src095 <= 32'hffffffff;
      src096 <= 31'h7fffffff;
      src097 <= 30'h3fffffff;
      src098 <= 29'h1fffffff;
      src099 <= 28'hfffffff;
      src100 <= 27'h7ffffff;
      src101 <= 26'h3ffffff;
      src102 <= 25'h1ffffff;
      src103 <= 24'hffffff;
      src104 <= 23'h7fffff;
      src105 <= 22'h3fffff;
      src106 <= 21'h1fffff;
      src107 <= 20'hfffff;
      src108 <= 19'h7ffff;
      src109 <= 18'h3ffff;
      src110 <= 17'h1ffff;
      src111 <= 16'hffff;
      src112 <= 15'h7fff;
      src113 <= 14'h3fff;
      src114 <= 13'h1fff;
      src115 <= 12'hfff;
      src116 <= 11'h7ff;
      src117 <= 10'h3ff;
      src118 <= 9'h1ff;
      src119 <= 8'hff;
      src120 <= 7'h7f;
      src121 <= 6'h3f;
      src122 <= 5'h1f;
      src123 <= 4'hf;
      src124 <= 3'h7;
      src125 <= 2'h3;
      src126 <= 1'h1;
      #1
      src000 <= 1'h1;
      src001 <= 2'h3;
      src002 <= 3'h0;
      src003 <= 4'h8;
      src004 <= 5'h1f;
      src005 <= 6'h33;
      src006 <= 7'h4d;
      src007 <= 8'hf4;
      src008 <= 9'h16e;
      src009 <= 10'h1bf;
      src010 <= 11'h23a;
      src011 <= 12'h904;
      src012 <= 13'h8f1;
      src013 <= 14'hc23;
      src014 <= 15'h4021;
      src015 <= 16'h4b3e;
      src016 <= 17'h13d97;
      src017 <= 18'hca44;
      src018 <= 19'h12e0c;
      src019 <= 20'ha90f9;
      src020 <= 21'h1e3796;
      src021 <= 22'hce3c6;
      src022 <= 23'h5a9211;
      src023 <= 24'hde4bc5;
      src024 <= 25'h143c911;
      src025 <= 26'h1a2c53a;
      src026 <= 27'h7a1d500;
      src027 <= 28'he2a8b42;
      src028 <= 29'h10abe7f0;
      src029 <= 30'h7f8c701;
      src030 <= 31'h3983ca8;
      src031 <= 32'hd71037d1;
      src032 <= 33'ha0116be5;
      src033 <= 34'h39ca5499d;
      src034 <= 35'h355485822;
      src035 <= 36'habaf3897a;
      src036 <= 37'hc101fbccc;
      src037 <= 38'h1e38c1962e;
      src038 <= 39'h728b0163c1;
      src039 <= 40'h291759edc3;
      src040 <= 41'h147fe43c49e;
      src041 <= 42'hdf7d41e602;
      src042 <= 43'h71e49a3e80e;
      src043 <= 44'hc51cc457821;
      src044 <= 45'h12943dfabc08;
      src045 <= 46'h183d2f120554;
      src046 <= 47'h2fcdd24bace4;
      src047 <= 48'hf3fb42930b33;
      src048 <= 49'h5bfa11af923d;
      src049 <= 50'h3215faef9c00b;
      src050 <= 51'h468ff864a7a50;
      src051 <= 52'he6b0346743741;
      src052 <= 53'h545995b7c709a;
      src053 <= 54'h3e43cd1d878f9f;
      src054 <= 55'h3e379530bcab0e;
      src055 <= 56'h3bf9064562be7f;
      src056 <= 57'he1c068b490b608;
      src057 <= 58'h2a908b62ba4b180;
      src058 <= 59'h19c16a00febd845;
      src059 <= 60'h4aef7ffc87a7463;
      src060 <= 61'h2e51d6c38018b47;
      src061 <= 62'h36accf412f175ff;
      src062 <= 63'h64264cd51ea45cd6;
      src063 <= 64'h1db53334fb0323a1;
      src064 <= 63'h589f8779b025244;
      src065 <= 62'h17ad2915f87f43fd;
      src066 <= 61'h7ede5feb7d6467b;
      src067 <= 60'h6bd0af37aaf0e89;
      src068 <= 59'h5d5143ade9b2b4;
      src069 <= 58'h367aad88b53031d;
      src070 <= 57'h67efac9edfa3da;
      src071 <= 56'h851438d5fdb76a;
      src072 <= 55'h38884411ebcd49;
      src073 <= 54'h2cd66e4d125e7f;
      src074 <= 53'hb8a546fa231e9;
      src075 <= 52'h142977795e986;
      src076 <= 51'h19d5f98b33c6e;
      src077 <= 50'h19847642aad48;
      src078 <= 49'h16f29429817c5;
      src079 <= 48'h56be91dc59ef;
      src080 <= 47'hedcc470f0e7;
      src081 <= 46'h2bd02975d279;
      src082 <= 45'h100b878b9f6b;
      src083 <= 44'he27ebe21368;
      src084 <= 43'h2ccaa6524ab;
      src085 <= 42'h3c50361524c;
      src086 <= 41'h1a3ae68690a;
      src087 <= 40'h9feae2025e;
      src088 <= 39'h5ba6208143;
      src089 <= 38'h20a859890c;
      src090 <= 37'hb0d9c2aa;
      src091 <= 36'ha143e2e04;
      src092 <= 35'hbd30291a;
      src093 <= 34'h28b5885ca;
      src094 <= 33'h2284b7a4;
      src095 <= 32'h7b59051b;
      src096 <= 31'h49b25ded;
      src097 <= 30'h2dfa4e02;
      src098 <= 29'h8785425;
      src099 <= 28'h9edf530;
      src100 <= 27'h635518f;
      src101 <= 26'h350ba60;
      src102 <= 25'h52a914;
      src103 <= 24'hc7c8;
      src104 <= 23'h313b32;
      src105 <= 22'h2acdac;
      src106 <= 21'ha3ebf;
      src107 <= 20'h7a94b;
      src108 <= 19'h391cf;
      src109 <= 18'h395c7;
      src110 <= 17'h183bc;
      src111 <= 16'hd42d;
      src112 <= 15'h813;
      src113 <= 14'h337d;
      src114 <= 13'h1ac4;
      src115 <= 12'h17f;
      src116 <= 11'h2a6;
      src117 <= 10'h390;
      src118 <= 9'h41;
      src119 <= 8'h84;
      src120 <= 7'h28;
      src121 <= 6'h39;
      src122 <= 5'h1f;
      src123 <= 4'h0;
      src124 <= 3'h0;
      src125 <= 2'h3;
      src126 <= 1'h1;
      #1
      src000 <= 1'h1;
      src001 <= 2'h3;
      src002 <= 3'h0;
      src003 <= 4'hd;
      src004 <= 5'hc;
      src005 <= 6'ha;
      src006 <= 7'h21;
      src007 <= 8'h7;
      src008 <= 9'h19b;
      src009 <= 10'h357;
      src010 <= 11'h50f;
      src011 <= 12'h1b;
      src012 <= 13'hdaa;
      src013 <= 14'h1d4;
      src014 <= 15'h9a;
      src015 <= 16'h3210;
      src016 <= 17'hc307;
      src017 <= 18'hf383;
      src018 <= 19'h32d1f;
      src019 <= 20'h9ad64;
      src020 <= 21'h11eb3c;
      src021 <= 22'h175305;
      src022 <= 23'h19a571;
      src023 <= 24'hf3828f;
      src024 <= 25'h1963785;
      src025 <= 26'ha6986d;
      src026 <= 27'h597aab;
      src027 <= 28'h8ca74ac;
      src028 <= 29'h1cfd9836;
      src029 <= 30'hed1dbf1;
      src030 <= 31'h41a93f90;
      src031 <= 32'h58d87776;
      src032 <= 33'hdf3277fd;
      src033 <= 34'h4c14982;
      src034 <= 35'h30a68e88e;
      src035 <= 36'h8ae55cdff;
      src036 <= 37'h148ef066d4;
      src037 <= 38'h2ef24dfdd8;
      src038 <= 39'h7ea7c5cb87;
      src039 <= 40'heae7180322;
      src040 <= 41'h1bda3e04b3b;
      src041 <= 42'h16d89b5b368;
      src042 <= 43'h60235354579;
      src043 <= 44'h950964ddb77;
      src044 <= 45'h8dc0247145f;
      src045 <= 46'h22bc26a97465;
      src046 <= 47'h5667555a4085;
      src047 <= 48'hbc01ca24be4d;
      src048 <= 49'h5ff4b7ef941c;
      src049 <= 50'h490a9edb95f2;
      src050 <= 51'h4505f0a8c46c7;
      src051 <= 52'h4c80429f2c3c7;
      src052 <= 53'h1719184a1eb1b7;
      src053 <= 54'h1098138c69778f;
      src054 <= 55'h1d69d94b1cb8bd;
      src055 <= 56'h9da26a0c5a876f;
      src056 <= 57'h135ef4c122411e6;
      src057 <= 58'h264d0575419eefc;
      src058 <= 59'h1bd09446a2b3200;
      src059 <= 60'hf65c370e89dc815;
      src060 <= 61'h1592ba4279585e69;
      src061 <= 62'hfe9e00b57f98d1e;
      src062 <= 63'h1db2b4527aa56a18;
      src063 <= 64'h7f6b8793b318ad4c;
      src064 <= 63'h4d4985dc09aedbd0;
      src065 <= 62'h3012b8cc90823eda;
      src066 <= 61'h436a2a516408169;
      src067 <= 60'h2b59cf4ceca2ee3;
      src068 <= 59'hfa7ee038974df5;
      src069 <= 58'h10143062830869;
      src070 <= 57'h1934264191b8adf;
      src071 <= 56'he5a7984a31b243;
      src072 <= 55'h7d161feb8f2056;
      src073 <= 54'h36261c379deda1;
      src074 <= 53'h1792be156af458;
      src075 <= 52'h8596dffc573d5;
      src076 <= 51'h6e6482aa50f4e;
      src077 <= 50'h2de3f31234efe;
      src078 <= 49'h41631d7173e5;
      src079 <= 48'he739869bdbd2;
      src080 <= 47'h1e7033a1d1c2;
      src081 <= 46'h32f07f411fed;
      src082 <= 45'hd4341a8a6e1;
      src083 <= 44'h158a41865bf;
      src084 <= 43'h374cc249558;
      src085 <= 42'h12b9f982188;
      src086 <= 41'hca1ac902ee;
      src087 <= 40'hc1755a3ac1;
      src088 <= 39'h26d3b564b0;
      src089 <= 38'h127ce71b48;
      src090 <= 37'h19905c053b;
      src091 <= 36'hf856f3d95;
      src092 <= 35'h5e345ac72;
      src093 <= 34'h3d5627386;
      src094 <= 33'h1ff88ec82;
      src095 <= 32'hdfec4623;
      src096 <= 31'h38018399;
      src097 <= 30'h13e009f;
      src098 <= 29'h15c62b68;
      src099 <= 28'ha2f2e6a;
      src100 <= 27'h52631db;
      src101 <= 26'h48a395;
      src102 <= 25'h97ed7c;
      src103 <= 24'h838606;
      src104 <= 23'h27e969;
      src105 <= 22'h30833d;
      src106 <= 21'h12d729;
      src107 <= 20'hf0dc6;
      src108 <= 19'h10fce;
      src109 <= 18'had59;
      src110 <= 17'h285c;
      src111 <= 16'h21f9;
      src112 <= 15'h399f;
      src113 <= 14'h10b4;
      src114 <= 13'h299;
      src115 <= 12'h99d;
      src116 <= 11'h3e;
      src117 <= 10'h396;
      src118 <= 9'h152;
      src119 <= 8'h52;
      src120 <= 7'h26;
      src121 <= 6'h3a;
      src122 <= 5'h17;
      src123 <= 4'hc;
      src124 <= 3'h0;
      src125 <= 2'h0;
      src126 <= 1'h0;
      #1
      src000 <= 1'h1;
      src001 <= 2'h1;
      src002 <= 3'h4;
      src003 <= 4'hd;
      src004 <= 5'h1e;
      src005 <= 6'h31;
      src006 <= 7'h3b;
      src007 <= 8'ha;
      src008 <= 9'h0;
      src009 <= 10'h174;
      src010 <= 11'h4d6;
      src011 <= 12'h824;
      src012 <= 13'h154a;
      src013 <= 14'h866;
      src014 <= 15'h7e56;
      src015 <= 16'h8625;
      src016 <= 17'h13612;
      src017 <= 18'h343bb;
      src018 <= 19'h62584;
      src019 <= 20'hc471a;
      src020 <= 21'h3fc0c;
      src021 <= 22'h14f73f;
      src022 <= 23'h209818;
      src023 <= 24'h7a57e0;
      src024 <= 25'h125fa7c;
      src025 <= 26'h2ac151d;
      src026 <= 27'he37052;
      src027 <= 28'h1265eb6;
      src028 <= 29'h1ece1e16;
      src029 <= 30'h357ca270;
      src030 <= 31'h2412579d;
      src031 <= 32'hb799ae8e;
      src032 <= 33'h1fc98c279;
      src033 <= 34'h69407be7;
      src034 <= 35'h79c9d03f3;
      src035 <= 36'he62fda854;
      src036 <= 37'h60c0a5967;
      src037 <= 38'h226c00984;
      src038 <= 39'h219e0df45b;
      src039 <= 40'ha5a1457899;
      src040 <= 41'hc758bf3b9e;
      src041 <= 42'he37d859725;
      src042 <= 43'hf6e19b5837;
      src043 <= 44'h97b9f3dd894;
      src044 <= 45'h18cfe96aa1af;
      src045 <= 46'h259bcca1a034;
      src046 <= 47'h1f1ecf6c9992;
      src047 <= 48'h138c306aa871;
      src048 <= 49'h1916fc838a145;
      src049 <= 50'h2f8ff71cff814;
      src050 <= 51'h30c32c1b199c4;
      src051 <= 52'hb68e37499b28c;
      src052 <= 53'h28f0bef2d9a38;
      src053 <= 54'h20b07f7c7550f2;
      src054 <= 55'h6d2ede6ac9d8a;
      src055 <= 56'h75955f374a6cc9;
      src056 <= 57'h952fde1d0ab994;
      src057 <= 58'h3605f2a90e639e1;
      src058 <= 59'h15831feec41e6f6;
      src059 <= 60'h35a3b55ef8d9ff0;
      src060 <= 61'h406ed7e6a677623;
      src061 <= 62'h352402a11965e435;
      src062 <= 63'h27f9e728c618fc1e;
      src063 <= 64'hf45da406bbf9bb01;
      src064 <= 63'h725c2675ca9571e4;
      src065 <= 62'h3db70476ac1ca75;
      src066 <= 61'h506c68640a978bf;
      src067 <= 60'h24023955a3da367;
      src068 <= 59'h5bf80671f12a0e9;
      src069 <= 58'h3c2a46b1182d23;
      src070 <= 57'h1643a0f586f1721;
      src071 <= 56'h51a082d8b5b41;
      src072 <= 55'h120d715da53b38;
      src073 <= 54'h1a9f0624aeba79;
      src074 <= 53'hd1b4a00d3d1af;
      src075 <= 52'h3f128e6a1a40b;
      src076 <= 51'h1d6dbf7b68ae;
      src077 <= 50'h2f3fa4b1347f6;
      src078 <= 49'h193db080e003;
      src079 <= 48'h5fbd2452bc39;
      src080 <= 47'h1cc5743c7e9d;
      src081 <= 46'h2c167a089ca8;
      src082 <= 45'h854421aa15e;
      src083 <= 44'hb9735475c5e;
      src084 <= 43'h79255c36c3d;
      src085 <= 42'h257f5fe0213;
      src086 <= 41'hbc53b53b92;
      src087 <= 40'h3414afe646;
      src088 <= 39'h284ec985ff;
      src089 <= 38'h28390a9016;
      src090 <= 37'hf82221345;
      src091 <= 36'h92f16fb50;
      src092 <= 35'h65f59aa2c;
      src093 <= 34'ha9c72e7b;
      src094 <= 33'hdc68d4fd;
      src095 <= 32'h99e8c828;
      src096 <= 31'h64d02759;
      src097 <= 30'h9f951be;
      src098 <= 29'h4af7dd7;
      src099 <= 28'h4398296;
      src100 <= 27'h6b944e0;
      src101 <= 26'h26524d5;
      src102 <= 25'h1aac055;
      src103 <= 24'h48d961;
      src104 <= 23'h6c148f;
      src105 <= 22'h2625c8;
      src106 <= 21'h16b12d;
      src107 <= 20'h2b4ae;
      src108 <= 19'h3f80c;
      src109 <= 18'h38ef9;
      src110 <= 17'h17a1e;
      src111 <= 16'h1d9f;
      src112 <= 15'h605d;
      src113 <= 14'h344d;
      src114 <= 13'h8a;
      src115 <= 12'hd59;
      src116 <= 11'h521;
      src117 <= 10'h387;
      src118 <= 9'hd0;
      src119 <= 8'hbe;
      src120 <= 7'h4b;
      src121 <= 6'h3c;
      src122 <= 5'h5;
      src123 <= 4'h5;
      src124 <= 3'h1;
      src125 <= 2'h2;
      src126 <= 1'h0;
      #1
      src000 <= 1'h0;
      src001 <= 2'h3;
      src002 <= 3'h6;
      src003 <= 4'h5;
      src004 <= 5'h1a;
      src005 <= 6'h37;
      src006 <= 7'h2c;
      src007 <= 8'h7e;
      src008 <= 9'h1d0;
      src009 <= 10'h2b9;
      src010 <= 11'h247;
      src011 <= 12'hb5f;
      src012 <= 13'h1d98;
      src013 <= 14'hb12;
      src014 <= 15'h7bb8;
      src015 <= 16'h6843;
      src016 <= 17'h12dcd;
      src017 <= 18'h3c6;
      src018 <= 19'h72f77;
      src019 <= 20'hec8ca;
      src020 <= 21'h7f69;
      src021 <= 22'h1bff7b;
      src022 <= 23'h4c6e6f;
      src023 <= 24'h3a9a23;
      src024 <= 25'h1346304;
      src025 <= 26'h13ff0da;
      src026 <= 27'h6c98f73;
      src027 <= 28'hf15feb1;
      src028 <= 29'h5ec639b;
      src029 <= 30'h3fb3f70d;
      src030 <= 31'h3b7c1f9a;
      src031 <= 32'h67c21355;
      src032 <= 33'h588d91d;
      src033 <= 34'hab2212c9;
      src034 <= 35'h400109824;
      src035 <= 36'hcb5c03f6f;
      src036 <= 37'h671d04b0f;
      src037 <= 38'h20bf1df687;
      src038 <= 39'h485a9414b8;
      src039 <= 40'h1215d38ca9;
      src040 <= 41'h1384332559d;
      src041 <= 42'h2b8889c8ae2;
      src042 <= 43'h3fcdc0520a4;
      src043 <= 44'h53bc31277fd;
      src044 <= 45'h1a8c116e8a64;
      src045 <= 46'h2514dc66a27b;
      src046 <= 47'h692a1af55c26;
      src047 <= 48'hce8c8b279c29;
      src048 <= 49'h12b4447534952;
      src049 <= 50'h2f974713eceb1;
      src050 <= 51'h2835b2347b24f;
      src051 <= 52'hc34a71eda4209;
      src052 <= 53'h8ee1c77cb1a27;
      src053 <= 54'h2d51c44c88b9d8;
      src054 <= 55'h79009ca1d20ebc;
      src055 <= 56'hd488f5be0a5a56;
      src056 <= 57'h1e8280a37cf8025;
      src057 <= 58'h28bc1818066b49b;
      src058 <= 59'hf6ab75f55b2e5c;
      src059 <= 60'h99b1de471a8c9c6;
      src060 <= 61'h35a9e2c7eda9ab9;
      src061 <= 62'h3451e1c3739076a;
      src062 <= 63'h78b61daf5afb9565;
      src063 <= 64'h65264961ab4414ae;
      src064 <= 63'ha8aa1e45c7cbc62;
      src065 <= 62'h1d041490e695f8ba;
      src066 <= 61'h126d593e92a651d7;
      src067 <= 60'h35fee3530f2c485;
      src068 <= 59'h75fd3536f1bdd07;
      src069 <= 58'h2a43daeb7626f49;
      src070 <= 57'hac4b2462565a95;
      src071 <= 56'hd7ea5b54a8762b;
      src072 <= 55'h6f6ddfaffe2554;
      src073 <= 54'h3940dc25e4979d;
      src074 <= 53'h8453050ea1324;
      src075 <= 52'he36442fd3b9f2;
      src076 <= 51'h638d5fbc59e92;
      src077 <= 50'h31dc57df0fe6b;
      src078 <= 49'he171bad3116b;
      src079 <= 48'h6473cbab5b51;
      src080 <= 47'hcbfb5c25d42;
      src081 <= 46'h31b5e7e3f52c;
      src082 <= 45'hefa0884fd16;
      src083 <= 44'h2b5a217cf25;
      src084 <= 43'h2fcdefa7864;
      src085 <= 42'h745d158e44;
      src086 <= 41'hb1ad7027cf;
      src087 <= 40'h91c061c99b;
      src088 <= 39'h5ae2091f49;
      src089 <= 38'h3a6953a115;
      src090 <= 37'h1f7460d20d;
      src091 <= 36'h679c45c38;
      src092 <= 35'h456525ce0;
      src093 <= 34'hacfeba4;
      src094 <= 33'hd742256;
      src095 <= 32'h598ca3b4;
      src096 <= 31'h4a30f7cd;
      src097 <= 30'he9a348;
      src098 <= 29'h8fc6d9f;
      src099 <= 28'h209bfec;
      src100 <= 27'h6d80ab0;
      src101 <= 26'h1c6ff3b;
      src102 <= 25'h19607e4;
      src103 <= 24'h71235d;
      src104 <= 23'h7425f4;
      src105 <= 22'h18af40;
      src106 <= 21'h15ba6d;
      src107 <= 20'h3465c;
      src108 <= 19'h15eb3;
      src109 <= 18'h28d5f;
      src110 <= 17'h14aad;
      src111 <= 16'he957;
      src112 <= 15'h533c;
      src113 <= 14'h20b4;
      src114 <= 13'h1d8;
      src115 <= 12'h16b;
      src116 <= 11'h30a;
      src117 <= 10'h2f3;
      src118 <= 9'h52;
      src119 <= 8'h6b;
      src120 <= 7'h58;
      src121 <= 6'h18;
      src122 <= 5'hc;
      src123 <= 4'h8;
      src124 <= 3'h4;
      src125 <= 2'h2;
      src126 <= 1'h1;
      #1
      src000 <= 1'h1;
      src001 <= 2'h3;
      src002 <= 3'h5;
      src003 <= 4'h7;
      src004 <= 5'h2;
      src005 <= 6'h27;
      src006 <= 7'h12;
      src007 <= 8'h4;
      src008 <= 9'h1d7;
      src009 <= 10'h3f6;
      src010 <= 11'h702;
      src011 <= 12'h184;
      src012 <= 13'h1a60;
      src013 <= 14'h3f2d;
      src014 <= 15'h75e4;
      src015 <= 16'he155;
      src016 <= 17'h78f5;
      src017 <= 18'haf57;
      src018 <= 19'h14dba;
      src019 <= 20'h7b774;
      src020 <= 21'h65199;
      src021 <= 22'h13af93;
      src022 <= 23'h69fcbe;
      src023 <= 24'h6d4b7c;
      src024 <= 25'h1c33712;
      src025 <= 26'h9dfd4f;
      src026 <= 27'h6d4ba69;
      src027 <= 28'hc9f81b7;
      src028 <= 29'h284bcec;
      src029 <= 30'h1716ffef;
      src030 <= 31'h3fee2fc7;
      src031 <= 32'h7d718591;
      src032 <= 33'h1deffed7a;
      src033 <= 34'h2ef38d426;
      src034 <= 35'h16f51ea78;
      src035 <= 36'he9acba588;
      src036 <= 37'h1142d01ba3;
      src037 <= 38'h23b56735e;
      src038 <= 39'h2c19518f87;
      src039 <= 40'hd4bb9e5a02;
      src040 <= 41'hdf3fafa217;
      src041 <= 42'hda8dce886;
      src042 <= 43'h6da83e9973b;
      src043 <= 44'h197dbedb42e;
      src044 <= 45'h189e1f2de275;
      src045 <= 46'h22e0a52ba0ce;
      src046 <= 47'h3ac45be12d09;
      src047 <= 48'h9078a91da2cd;
      src048 <= 49'h42573d798f0b;
      src049 <= 50'h275cc84a5b1c3;
      src050 <= 51'h53ca8acb5959f;
      src051 <= 52'hbf13a3bcd6aec;
      src052 <= 53'h1ebcbda0e624f1;
      src053 <= 54'h1192a62bdfb727;
      src054 <= 55'h3f7bacf4bb315;
      src055 <= 56'hbbe5c053f04099;
      src056 <= 57'h9ef80e6544c97d;
      src057 <= 58'h16a03b5f9cb2ee8;
      src058 <= 59'h22b56be1392a255;
      src059 <= 60'h69baec4c3d9b3b0;
      src060 <= 61'h1fca8b99c6596f7f;
      src061 <= 62'h1e1ed48836a52df9;
      src062 <= 63'h21d32e24bb891746;
      src063 <= 64'h7d3c279b5bce228b;
      src064 <= 63'h33c14694f06ea18;
      src065 <= 62'h1c2b5f18f568c9c6;
      src066 <= 61'h1fa925bde10b4aad;
      src067 <= 60'hf63a809bcc4616d;
      src068 <= 59'h505e9c98bc88bcf;
      src069 <= 58'h212c196142a6c95;
      src070 <= 57'h1894f7f4aaeb212;
      src071 <= 56'h1e4ce1f19b43da;
      src072 <= 55'h9cd3b356af737;
      src073 <= 54'h2becd73fe65f90;
      src074 <= 53'h1c3c8adceb2013;
      src075 <= 52'h852cb39d5b552;
      src076 <= 51'h4e0e1298e9a79;
      src077 <= 50'h2d9d2045892c1;
      src078 <= 49'h9ad8a1645f58;
      src079 <= 48'hb415a79b46a;
      src080 <= 47'h6490fb2de1e;
      src081 <= 46'h5c13dd0c866;
      src082 <= 45'he73032f594d;
      src083 <= 44'h22153a081a6;
      src084 <= 43'hffd22a3a62;
      src085 <= 42'h361a9fa4ea6;
      src086 <= 41'hddec071cf1;
      src087 <= 40'hde72ef7dce;
      src088 <= 39'h5b245db6ca;
      src089 <= 38'h164fdc1351;
      src090 <= 37'h15a629d332;
      src091 <= 36'hc689c0559;
      src092 <= 35'h6027752fe;
      src093 <= 34'h2e413961f;
      src094 <= 33'h1b476998d;
      src095 <= 32'hc2537638;
      src096 <= 31'h1f626a97;
      src097 <= 30'h3457f15c;
      src098 <= 29'h18faa81f;
      src099 <= 28'h57b6ae4;
      src100 <= 27'hcbd31;
      src101 <= 26'h11b16de;
      src102 <= 25'h97b952;
      src103 <= 24'h28c78b;
      src104 <= 23'h547e39;
      src105 <= 22'h1e627b;
      src106 <= 21'hb4812;
      src107 <= 20'h7e5bd;
      src108 <= 19'h5a02;
      src109 <= 18'h159ca;
      src110 <= 17'hac5a;
      src111 <= 16'h282f;
      src112 <= 15'h6d5b;
      src113 <= 14'hd44;
      src114 <= 13'h1d47;
      src115 <= 12'h4cd;
      src116 <= 11'ha4;
      src117 <= 10'h205;
      src118 <= 9'h15c;
      src119 <= 8'hc0;
      src120 <= 7'h6;
      src121 <= 6'h4;
      src122 <= 5'h1f;
      src123 <= 4'h2;
      src124 <= 3'h5;
      src125 <= 2'h2;
      src126 <= 1'h0;
      #1
      src000 <= 1'h1;
      src001 <= 2'h1;
      src002 <= 3'h5;
      src003 <= 4'h5;
      src004 <= 5'h19;
      src005 <= 6'h2b;
      src006 <= 7'h45;
      src007 <= 8'hfc;
      src008 <= 9'h192;
      src009 <= 10'h1e;
      src010 <= 11'h4f8;
      src011 <= 12'h939;
      src012 <= 13'h1e02;
      src013 <= 14'h478;
      src014 <= 15'h432f;
      src015 <= 16'h139c;
      src016 <= 17'h1d2dc;
      src017 <= 18'h32917;
      src018 <= 19'h1eb95;
      src019 <= 20'hcebc1;
      src020 <= 21'h162e82;
      src021 <= 22'h3f7d17;
      src022 <= 23'hd1853;
      src023 <= 24'ha9710;
      src024 <= 25'h1179a56;
      src025 <= 26'h463135;
      src026 <= 27'h4100e66;
      src027 <= 28'h945dba8;
      src028 <= 29'hd4117dd;
      src029 <= 30'h2b8e4ebc;
      src030 <= 31'h62d59938;
      src031 <= 32'hf8cc3f3b;
      src032 <= 33'h357f0a64;
      src033 <= 34'h1ecadbb86;
      src034 <= 35'h25a7583c0;
      src035 <= 36'h4e642965c;
      src036 <= 37'h3d0fce922;
      src037 <= 38'h13909b471c;
      src038 <= 39'h58f3ca5f64;
      src039 <= 40'h955cfa38b1;
      src040 <= 41'h12ca02ebb76;
      src041 <= 42'h3f552b04994;
      src042 <= 43'h675c8649f78;
      src043 <= 44'hdca99c7abea;
      src044 <= 45'hae1fccae6b8;
      src045 <= 46'h388f0b2975c6;
      src046 <= 47'h576220379089;
      src047 <= 48'h4c5edec31ef;
      src048 <= 49'h107c8c7537df5;
      src049 <= 50'h8fdd300a2187;
      src050 <= 51'h475956c835975;
      src051 <= 52'h206722b7bde99;
      src052 <= 53'h189ee79ae445e0;
      src053 <= 54'h37a234c1378e75;
      src054 <= 55'h4fb7c34408c04c;
      src055 <= 56'h6fb2e48f3531c;
      src056 <= 57'h11f2bddb7c97da8;
      src057 <= 58'h210c651f23db306;
      src058 <= 59'h5163de18df7a267;
      src059 <= 60'haf3d348fd768f63;
      src060 <= 61'h1ba0e9ecc857d8c3;
      src061 <= 62'h12237677caa0a679;
      src062 <= 63'h1847803d840fccb;
      src063 <= 64'h82e7448cc0037457;
      src064 <= 63'h5c66a9bb62574c5a;
      src065 <= 62'h34b08056e994f3e6;
      src066 <= 61'he9c805fc29ed120;
      src067 <= 60'h808c98e65a3ae4;
      src068 <= 59'h7f3ab7db3390a6e;
      src069 <= 58'h1fe59a7bc39e1b3;
      src070 <= 57'h1190f5c3df8eeef;
      src071 <= 56'h27e5b96b83f00f;
      src072 <= 55'h72bbe792b95731;
      src073 <= 54'h398e43b6bca2a2;
      src074 <= 53'ha86f030331476;
      src075 <= 52'h816004598244b;
      src076 <= 51'h1733753e83663;
      src077 <= 50'h3db74e98ce25;
      src078 <= 49'hb3b7e15aa2c;
      src079 <= 48'h8049c334f558;
      src080 <= 47'h62f965dcac6c;
      src081 <= 46'h31d3ac4ebce0;
      src082 <= 45'h275d2928f4b;
      src083 <= 44'hee3952b1ee1;
      src084 <= 43'h207919c21ed;
      src085 <= 42'h29f4741ee56;
      src086 <= 41'h18d26eeeba;
      src087 <= 40'hf265e96753;
      src088 <= 39'ha22a5a421;
      src089 <= 38'h2cdd6d47e4;
      src090 <= 37'h5c6be596;
      src091 <= 36'h611c272d8;
      src092 <= 35'h1b7a02afd;
      src093 <= 34'h789a2829;
      src094 <= 33'h1067fece7;
      src095 <= 32'ha2b4d215;
      src096 <= 31'h680aee2a;
      src097 <= 30'h1231613a;
      src098 <= 29'h97077d9;
      src099 <= 28'hcef3bc1;
      src100 <= 27'h4e5c6dd;
      src101 <= 26'h7a91b0;
      src102 <= 25'ha6d259;
      src103 <= 24'h403221;
      src104 <= 23'h224af3;
      src105 <= 22'h3d8de5;
      src106 <= 21'h2fd5b;
      src107 <= 20'h1641d;
      src108 <= 19'h6323c;
      src109 <= 18'h17117;
      src110 <= 17'h160f8;
      src111 <= 16'h2a64;
      src112 <= 15'h14aa;
      src113 <= 14'h1653;
      src114 <= 13'h10ff;
      src115 <= 12'h673;
      src116 <= 11'h42c;
      src117 <= 10'h29f;
      src118 <= 9'h103;
      src119 <= 8'h84;
      src120 <= 7'h74;
      src121 <= 6'h13;
      src122 <= 5'h1c;
      src123 <= 4'h4;
      src124 <= 3'h0;
      src125 <= 2'h1;
      src126 <= 1'h0;
      #1
      src000 <= 1'h1;
      src001 <= 2'h0;
      src002 <= 3'h3;
      src003 <= 4'he;
      src004 <= 5'hf;
      src005 <= 6'h3a;
      src006 <= 7'h28;
      src007 <= 8'haa;
      src008 <= 9'h8a;
      src009 <= 10'h3cf;
      src010 <= 11'hea;
      src011 <= 12'h2a3;
      src012 <= 13'h15f9;
      src013 <= 14'h50;
      src014 <= 15'h147a;
      src015 <= 16'h353d;
      src016 <= 17'h1b5ff;
      src017 <= 18'h2d18d;
      src018 <= 19'h739ac;
      src019 <= 20'habeef;
      src020 <= 21'h183239;
      src021 <= 22'h2e57d0;
      src022 <= 23'h1e6cbd;
      src023 <= 24'h45b002;
      src024 <= 25'h1447f36;
      src025 <= 26'h2e8ab5;
      src026 <= 27'h2ebed37;
      src027 <= 28'h400d183;
      src028 <= 29'h13a9607;
      src029 <= 30'h2b3ff62f;
      src030 <= 31'h317eeb1d;
      src031 <= 32'hb4cba0a;
      src032 <= 33'ha5387901;
      src033 <= 34'h2b2e74e77;
      src034 <= 35'h6cbf8e26a;
      src035 <= 36'h1e963544a;
      src036 <= 37'h162b0c9fdd;
      src037 <= 38'h9ed469bf4;
      src038 <= 39'hd688181a8;
      src039 <= 40'hb570d22718;
      src040 <= 41'h1a674219d3e;
      src041 <= 42'h3e2e402534;
      src042 <= 43'h30c439f4b86;
      src043 <= 44'hc67f30459cc;
      src044 <= 45'h16e3106861d3;
      src045 <= 46'hfca18a77594;
      src046 <= 47'h59cd06b42b6f;
      src047 <= 48'h5aab05765983;
      src048 <= 49'hdf9e5a1bdae;
      src049 <= 50'h3a6dc52a33c33;
      src050 <= 51'h7efbeb1e186d7;
      src051 <= 52'h2930c79fe0a1b;
      src052 <= 53'h34f71dba45b5e;
      src053 <= 54'h21912aeceb9505;
      src054 <= 55'h1880fa840fbb0b;
      src055 <= 56'haacf501480f037;
      src056 <= 57'h1e2b21c19365f61;
      src057 <= 58'h43b8fff7d870b6;
      src058 <= 59'h497e28ace03a34d;
      src059 <= 60'h12d7f5ff5b7751f;
      src060 <= 61'h181ba140002f9cc4;
      src061 <= 62'h141401b85672ebc7;
      src062 <= 63'h259a2b28b22b8974;
      src063 <= 64'hf212cc6f540988e7;
      src064 <= 63'h65ea29d1adae7e45;
      src065 <= 62'h1cfb836a0b4ea16d;
      src066 <= 61'h150746a04815642c;
      src067 <= 60'hb4441d63cf9d1fe;
      src068 <= 59'h29e316a39ddc477;
      src069 <= 58'h35db102e0db22d3;
      src070 <= 57'h174015c7680891b;
      src071 <= 56'hc5e4a52353d455;
      src072 <= 55'h29821003729e33;
      src073 <= 54'h1602dccd34bcd7;
      src074 <= 53'h9873bfff83cec;
      src075 <= 52'hce2904fe973d;
      src076 <= 51'h52c55d2f74429;
      src077 <= 50'h79282951fe0;
      src078 <= 49'h305609c64c1d;
      src079 <= 48'h4b9e9c899296;
      src080 <= 47'h2734c7405255;
      src081 <= 46'h359906c4e109;
      src082 <= 45'h174c2348e1b7;
      src083 <= 44'h6ee829fe7ba;
      src084 <= 43'h6678889832c;
      src085 <= 42'h10912b34a24;
      src086 <= 41'h167a89f5916;
      src087 <= 40'h31f74f1905;
      src088 <= 39'h3e6fa00319;
      src089 <= 38'h30789c3c72;
      src090 <= 37'hf65141471;
      src091 <= 36'hfa53011a2;
      src092 <= 35'h194d50a99;
      src093 <= 34'h2d5e8b89c;
      src094 <= 33'h1ff7acd86;
      src095 <= 32'h3cad275a;
      src096 <= 31'ha515e87;
      src097 <= 30'h292936a2;
      src098 <= 29'h190277cc;
      src099 <= 28'h369c285;
      src100 <= 27'hc78c2f;
      src101 <= 26'h127561f;
      src102 <= 25'h191d902;
      src103 <= 24'hdb82a;
      src104 <= 23'h6bc9e9;
      src105 <= 22'h32515e;
      src106 <= 21'h1bb58f;
      src107 <= 20'h35aac;
      src108 <= 19'h75ef8;
      src109 <= 18'h3b226;
      src110 <= 17'ha540;
      src111 <= 16'h56d6;
      src112 <= 15'h572a;
      src113 <= 14'h3cb7;
      src114 <= 13'h1a4f;
      src115 <= 12'h516;
      src116 <= 11'h48a;
      src117 <= 10'he6;
      src118 <= 9'h179;
      src119 <= 8'hb0;
      src120 <= 7'h24;
      src121 <= 6'h2d;
      src122 <= 5'h1e;
      src123 <= 4'h1;
      src124 <= 3'h3;
      src125 <= 2'h2;
      src126 <= 1'h0;
      #1
      src000 <= 1'h1;
      src001 <= 2'h2;
      src002 <= 3'h6;
      src003 <= 4'h1;
      src004 <= 5'h12;
      src005 <= 6'h37;
      src006 <= 7'h8;
      src007 <= 8'hd2;
      src008 <= 9'h113;
      src009 <= 10'h300;
      src010 <= 11'h354;
      src011 <= 12'hb19;
      src012 <= 13'h896;
      src013 <= 14'h10ea;
      src014 <= 15'h1c3c;
      src015 <= 16'hb6c3;
      src016 <= 17'ha9bc;
      src017 <= 18'h3ff3;
      src018 <= 19'h6e3a5;
      src019 <= 20'hcbfab;
      src020 <= 21'h1daa4c;
      src021 <= 22'h9bfe6;
      src022 <= 23'h13ec57;
      src023 <= 24'hd9d1af;
      src024 <= 25'h8d9eb6;
      src025 <= 26'h15a96d5;
      src026 <= 27'h2728ec9;
      src027 <= 28'h6a38b55;
      src028 <= 29'ha86b3a1;
      src029 <= 30'h1d374789;
      src030 <= 31'h79be4e5;
      src031 <= 32'h867a4ac9;
      src032 <= 33'h1d1a8d7b0;
      src033 <= 34'h2bc6284a8;
      src034 <= 35'h4dcfbde0a;
      src035 <= 36'h5e63317c3;
      src036 <= 37'h9b1f5d7d0;
      src037 <= 38'h30e983cc1d;
      src038 <= 39'h3c4e245cf7;
      src039 <= 40'hc1fe1c51e5;
      src040 <= 41'h18f58b5f052;
      src041 <= 42'h3c5f2ded00f;
      src042 <= 43'h4e682f4b48a;
      src043 <= 44'hd1ff6f25926;
      src044 <= 45'h1a00fef06b04;
      src045 <= 46'hc81d01cf935;
      src046 <= 47'h25cc276d7e19;
      src047 <= 48'h36b08461f840;
      src048 <= 49'h111141c769e1f;
      src049 <= 50'h1595e9d4319b5;
      src050 <= 51'h15db4603803f3;
      src051 <= 52'h12715cb18d6a4;
      src052 <= 53'h762b002af3382;
      src053 <= 54'h2e5b78e4751694;
      src054 <= 55'h517fa07b0f78c1;
      src055 <= 56'hbcf9f573df770a;
      src056 <= 57'hea3470c6962905;
      src057 <= 58'h145ba79ec3826bc;
      src058 <= 59'h6999e12b02237e;
      src059 <= 60'h5568cbdd97d2b38;
      src060 <= 61'h1a2b70a38463416a;
      src061 <= 62'h381675df3544f189;
      src062 <= 63'h439ddd7467af36d9;
      src063 <= 64'h96625aa1056b565f;
      src064 <= 63'h636241c3eb6ec9e0;
      src065 <= 62'hb1c192ecd6665d8;
      src066 <= 61'h1568e84a67ba6b1a;
      src067 <= 60'he93a8c0df983779;
      src068 <= 59'h7add8fe0a02da60;
      src069 <= 58'hd07f909eb88325;
      src070 <= 57'h1f60bf381eb88e5;
      src071 <= 56'hf202f364e322cf;
      src072 <= 55'h2e573843eb280e;
      src073 <= 54'h146bcc5d443821;
      src074 <= 53'h93160eab3c4d8;
      src075 <= 52'h233f874f8c57b;
      src076 <= 51'h1188af660ffd5;
      src077 <= 50'h3255d7a658abe;
      src078 <= 49'h10fe6179d221d;
      src079 <= 48'h75947b777bf2;
      src080 <= 47'h1c62d0813d92;
      src081 <= 46'h120e4bf41e10;
      src082 <= 45'h8df181a218e;
      src083 <= 44'h460aa61353a;
      src084 <= 43'h1c32d116fe;
      src085 <= 42'h3ec9a0a80be;
      src086 <= 41'h15fc7afae8f;
      src087 <= 40'h31df61c534;
      src088 <= 39'h1af8c96a9;
      src089 <= 38'h1d3ddf55b2;
      src090 <= 37'h13fbf70946;
      src091 <= 36'h74642cddb;
      src092 <= 35'h7024bfe48;
      src093 <= 34'h2ed3032ed;
      src094 <= 33'h17776c3a;
      src095 <= 32'h6c1b6811;
      src096 <= 31'h5e146c30;
      src097 <= 30'h30c9eda8;
      src098 <= 29'h94f7dcd;
      src099 <= 28'h76980e6;
      src100 <= 27'h49b3fe6;
      src101 <= 26'h19830b0;
      src102 <= 25'h1ecaa99;
      src103 <= 24'hb7e4dd;
      src104 <= 23'h486c0a;
      src105 <= 22'h31320c;
      src106 <= 21'h84795;
      src107 <= 20'h3d29d;
      src108 <= 19'h66b48;
      src109 <= 18'h2d729;
      src110 <= 17'h1e245;
      src111 <= 16'h7511;
      src112 <= 15'h5fba;
      src113 <= 14'h2deb;
      src114 <= 13'h1ba4;
      src115 <= 12'h8e0;
      src116 <= 11'h5bf;
      src117 <= 10'h334;
      src118 <= 9'h121;
      src119 <= 8'h35;
      src120 <= 7'h7a;
      src121 <= 6'h25;
      src122 <= 5'h7;
      src123 <= 4'he;
      src124 <= 3'h2;
      src125 <= 2'h2;
      src126 <= 1'h0;
      #1
      src000 <= 1'h0;
      src001 <= 2'h2;
      src002 <= 3'h7;
      src003 <= 4'h7;
      src004 <= 5'h7;
      src005 <= 6'h31;
      src006 <= 7'h63;
      src007 <= 8'hed;
      src008 <= 9'h1d8;
      src009 <= 10'h1c3;
      src010 <= 11'h663;
      src011 <= 12'h9f5;
      src012 <= 13'h1f25;
      src013 <= 14'h1dc7;
      src014 <= 15'h5084;
      src015 <= 16'hd7;
      src016 <= 17'h5e19;
      src017 <= 18'h3c62d;
      src018 <= 19'h51306;
      src019 <= 20'hc9dd8;
      src020 <= 21'he8d5d;
      src021 <= 22'h373684;
      src022 <= 23'hc72fe;
      src023 <= 24'h14b406;
      src024 <= 25'h1a04247;
      src025 <= 26'hbf717f;
      src026 <= 27'h437249f;
      src027 <= 28'h668def8;
      src028 <= 29'h14ea7b17;
      src029 <= 30'h16db6f10;
      src030 <= 31'h1cf4a8ed;
      src031 <= 32'hb2daa1f6;
      src032 <= 33'h73c36ba;
      src033 <= 34'hf3f05323;
      src034 <= 35'h60212585b;
      src035 <= 36'h88da091b;
      src036 <= 37'h7213124bd;
      src037 <= 38'h19e998952c;
      src038 <= 39'h327751b3fa;
      src039 <= 40'hd9073286;
      src040 <= 41'h446a4ace0e;
      src041 <= 42'h16a89745cd7;
      src042 <= 43'h3bfed0d0418;
      src043 <= 44'hc386a594b07;
      src044 <= 45'h1be400183cfe;
      src045 <= 46'h30cc35c9599f;
      src046 <= 47'h44f2f45c8840;
      src047 <= 48'h2f21845c21e7;
      src048 <= 49'h1176b1a7e256d;
      src049 <= 50'h3080122ca9fe8;
      src050 <= 51'h339fb51cd2c07;
      src051 <= 52'h3d9d6801841f4;
      src052 <= 53'h6c1028f41d3e4;
      src053 <= 54'hff12979801aaa;
      src054 <= 55'h7844c2729bd820;
      src055 <= 56'he8e8fe2dbdb6e5;
      src056 <= 57'h15bf88c8c3af69e;
      src057 <= 58'h35469f420fe652b;
      src058 <= 59'h60924d241229d75;
      src059 <= 60'habd2e31816480fa;
      src060 <= 61'hef2acfadcff697d;
      src061 <= 62'h1fcdde7e742c5905;
      src062 <= 63'h7b056d0259de5319;
      src063 <= 64'hef617cacc674d244;
      src064 <= 63'h726e8017061f5679;
      src065 <= 62'h1cab7dd472323dc9;
      src066 <= 61'hf6d84bd6df2fc82;
      src067 <= 60'hf457c0940d2d16f;
      src068 <= 59'h241813e799fde33;
      src069 <= 58'h386fb3d3a6f36fa;
      src070 <= 57'h1709dd84894d9fc;
      src071 <= 56'hf8ed4ba73e3f3b;
      src072 <= 55'h26184cedf6b1e0;
      src073 <= 54'h18037f166a1a98;
      src074 <= 53'h7db3bac546740;
      src075 <= 52'h1e34df239fbb0;
      src076 <= 51'h57c2727b51ee7;
      src077 <= 50'h2acef09642b31;
      src078 <= 49'ha434ce1f4081;
      src079 <= 48'hc7d577f63854;
      src080 <= 47'h3008ad830951;
      src081 <= 46'h3f8069560c06;
      src082 <= 45'hab8312a4c3c;
      src083 <= 44'h18264119d38;
      src084 <= 43'h56cf60ce881;
      src085 <= 42'h180855a7d8d;
      src086 <= 41'h14fb9534807;
      src087 <= 40'h4d6f1d5baf;
      src088 <= 39'h7e9e203161;
      src089 <= 38'h470fe3cfc;
      src090 <= 37'h1f3e332f35;
      src091 <= 36'had7f14ec2;
      src092 <= 35'h3246b7d9;
      src093 <= 34'hb2591c4;
      src094 <= 33'h2258edf3;
      src095 <= 32'haf3cb9d0;
      src096 <= 31'h6cef5e55;
      src097 <= 30'h24a881f6;
      src098 <= 29'h15a43dd3;
      src099 <= 28'hfca2d1b;
      src100 <= 27'h31307e4;
      src101 <= 26'h14e41b7;
      src102 <= 25'h17d94e0;
      src103 <= 24'hb68b9e;
      src104 <= 23'h702a5b;
      src105 <= 22'h320651;
      src106 <= 21'h1c16eb;
      src107 <= 20'ha292e;
      src108 <= 19'h77f45;
      src109 <= 18'h89e0;
      src110 <= 17'h961a;
      src111 <= 16'h7086;
      src112 <= 15'h1d01;
      src113 <= 14'h13f0;
      src114 <= 13'h1938;
      src115 <= 12'hed8;
      src116 <= 11'h35c;
      src117 <= 10'h2f1;
      src118 <= 9'h2f;
      src119 <= 8'ha;
      src120 <= 7'h67;
      src121 <= 6'h1a;
      src122 <= 5'h5;
      src123 <= 4'hd;
      src124 <= 3'h6;
      src125 <= 2'h1;
      src126 <= 1'h0;
      #1
      src000 <= 1'h0;
      src001 <= 2'h3;
      src002 <= 3'h4;
      src003 <= 4'hc;
      src004 <= 5'h4;
      src005 <= 6'ha;
      src006 <= 7'h7e;
      src007 <= 8'h7;
      src008 <= 9'hd0;
      src009 <= 10'h35a;
      src010 <= 11'h5c2;
      src011 <= 12'h9fc;
      src012 <= 13'h55b;
      src013 <= 14'h2f9;
      src014 <= 15'h3d37;
      src015 <= 16'he47;
      src016 <= 17'h17855;
      src017 <= 18'h13a1f;
      src018 <= 19'h773b8;
      src019 <= 20'h844c1;
      src020 <= 21'h70d47;
      src021 <= 22'h393c4e;
      src022 <= 23'h4748f7;
      src023 <= 24'h70660a;
      src024 <= 25'h187e710;
      src025 <= 26'h3128eba;
      src026 <= 27'h56fb5c7;
      src027 <= 28'h74e4973;
      src028 <= 29'h10e3722c;
      src029 <= 30'hb639aa5;
      src030 <= 31'hb44361f;
      src031 <= 32'h27a0008c;
      src032 <= 33'h19045a445;
      src033 <= 34'h37abc9f0b;
      src034 <= 35'h651c6a2e4;
      src035 <= 36'h30637fdca;
      src036 <= 37'h8f64e8f4a;
      src037 <= 38'h12c2fab184;
      src038 <= 39'h7e299cb48;
      src039 <= 40'h7e6e05724d;
      src040 <= 41'h10e45a16970;
      src041 <= 42'hec62614790;
      src042 <= 43'h4aa5804a881;
      src043 <= 44'h1e88abb572c;
      src044 <= 45'he48d5f52c0;
      src045 <= 46'h2101dcebef56;
      src046 <= 47'h233e54e27ea6;
      src047 <= 48'h32dafec24805;
      src048 <= 49'h1018f1152797e;
      src049 <= 50'hd561920c904e;
      src050 <= 51'h13389854ca896;
      src051 <= 52'h41ab8961139cf;
      src052 <= 53'h237da7c3ad037;
      src053 <= 54'h1c9818c82a6c15;
      src054 <= 55'h18c8ec58ea0417;
      src055 <= 56'h6f1612b5178761;
      src056 <= 57'hb57190fedcb8f9;
      src057 <= 58'h1d75adef63d307c;
      src058 <= 59'h338f4ac66270136;
      src059 <= 60'he0c28dfbecba4c8;
      src060 <= 61'ha1c0aec5931c9b4;
      src061 <= 62'h19b393aada2e6e6c;
      src062 <= 63'h773a13fb37503d77;
      src063 <= 64'h53fd2516d1bfbaba;
      src064 <= 63'h8fce7af52c1b3c7;
      src065 <= 62'h256d83cc039d60ba;
      src066 <= 61'h75691d3cda840fd;
      src067 <= 60'hb1540708dff06d2;
      src068 <= 59'h72f7892dd7516f5;
      src069 <= 58'h351232e16c2b4aa;
      src070 <= 57'h1a2fefdd4dc2301;
      src071 <= 56'h2926941f69cd43;
      src072 <= 55'h2c941552fa3935;
      src073 <= 54'h1eda654bebcf4f;
      src074 <= 53'h1bf717a0d9da58;
      src075 <= 52'h100c7496749fb;
      src076 <= 51'h44f06d87d3afc;
      src077 <= 50'h2890f5028361f;
      src078 <= 49'h319849954cf1;
      src079 <= 48'h47b084403b37;
      src080 <= 47'h6b29637c3644;
      src081 <= 46'h207139b66d71;
      src082 <= 45'h1404f367dbe2;
      src083 <= 44'hfa988653e42;
      src084 <= 43'h72ee3aeb12e;
      src085 <= 42'hfbb550f221;
      src086 <= 41'h17f6c749cf4;
      src087 <= 40'h760d20f686;
      src088 <= 39'h627a31a27c;
      src089 <= 38'h1e07d5e121;
      src090 <= 37'h1314c30b50;
      src091 <= 36'h700b1433;
      src092 <= 35'h169f5a741;
      src093 <= 34'h186ff76d1;
      src094 <= 33'h17ff5101d;
      src095 <= 32'h44bfc434;
      src096 <= 31'h6e771359;
      src097 <= 30'h3c40983e;
      src098 <= 29'h3bc16db;
      src099 <= 28'h5416408;
      src100 <= 27'h5b7801e;
      src101 <= 26'h19ea504;
      src102 <= 25'hff32cb;
      src103 <= 24'h4d6395;
      src104 <= 23'h38a7ac;
      src105 <= 22'h2681e5;
      src106 <= 21'h94c8f;
      src107 <= 20'h5f602;
      src108 <= 19'h401a2;
      src109 <= 18'h37cf;
      src110 <= 17'hb999;
      src111 <= 16'h771b;
      src112 <= 15'h6ad8;
      src113 <= 14'h1413;
      src114 <= 13'hf93;
      src115 <= 12'h41f;
      src116 <= 11'h2b0;
      src117 <= 10'h1fb;
      src118 <= 9'h132;
      src119 <= 8'ha;
      src120 <= 7'h75;
      src121 <= 6'h19;
      src122 <= 5'h3;
      src123 <= 4'hd;
      src124 <= 3'h2;
      src125 <= 2'h3;
      src126 <= 1'h1;
   end
endmodule

