module compressor(
      input wire [31:0] src00,
      input wire [31:0] src01,
      input wire [31:0] src02,
      input wire [31:0] src03,
      input wire [31:0] src04,
      input wire [31:0] src05,
      input wire [31:0] src06,
      input wire [31:0] src07,
      input wire [31:0] src08,
      input wire [31:0] src09,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      output wire [1:0] dst00,
      output wire [0:0] dst01,
      output wire [1:0] dst02,
      output wire [1:0] dst03,
      output wire [0:0] dst04,
      output wire [1:0] dst05,
      output wire [1:0] dst06,
      output wire [1:0] dst07,
      output wire [1:0] dst08,
      output wire [1:0] dst09,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [0:0] dst35,
      output wire [0:0] dst36
   );
   wire [51:0] stage00;
   wire [49:0] stage01;
   wire [56:0] stage02;
   wire [60:0] stage03;
   wire [70:0] stage04;
   wire [61:0] stage05;
   wire [51:0] stage06;
   wire [61:0] stage07;
   wire [56:0] stage08;
   wire [70:0] stage09;
   wire [62:0] stage10;
   wire [56:0] stage11;
   wire [57:0] stage12;
   wire [60:0] stage13;
   wire [59:0] stage14;
   wire [57:0] stage15;
   wire [66:0] stage16;
   wire [54:0] stage17;
   wire [57:0] stage18;
   wire [60:0] stage19;
   wire [58:0] stage20;
   wire [57:0] stage21;
   wire [60:0] stage22;
   wire [63:0] stage23;
   wire [62:0] stage24;
   wire [60:0] stage25;
   wire [67:0] stage26;
   wire [70:0] stage27;
   wire [66:0] stage28;
   wire [61:0] stage29;
   wire [66:0] stage30;
   wire [70:0] stage31;
   wire [17:0] stage32;
   wire [14:0] stage33;
   wire [4:0] stage34;
   wire [2:0] stage35;
   wire [0:0] stage36;
   assign stage00[31:0] = src00;
   assign stage01[31:0] = src01;
   assign stage02[31:0] = src02;
   assign stage03[31:0] = src03;
   assign stage04[31:0] = src04;
   assign stage05[31:0] = src05;
   assign stage06[31:0] = src06;
   assign stage07[31:0] = src07;
   assign stage08[31:0] = src08;
   assign stage09[31:0] = src09;
   assign stage10[31:0] = src10;
   assign stage11[31:0] = src11;
   assign stage12[31:0] = src12;
   assign stage13[31:0] = src13;
   assign stage14[31:0] = src14;
   assign stage15[31:0] = src15;
   assign stage16[31:0] = src16;
   assign stage17[31:0] = src17;
   assign stage18[31:0] = src18;
   assign stage19[31:0] = src19;
   assign stage20[31:0] = src20;
   assign stage21[31:0] = src21;
   assign stage22[31:0] = src22;
   assign stage23[31:0] = src23;
   assign stage24[31:0] = src24;
   assign stage25[31:0] = src25;
   assign stage26[31:0] = src26;
   assign stage27[31:0] = src27;
   assign stage28[31:0] = src28;
   assign stage29[31:0] = src29;
   assign stage30[31:0] = src30;
   assign stage31[31:0] = src31;
   assign dst00 = stage00[51:50];
   assign dst01 = stage01[49:49];
   assign dst02 = stage02[56:55];
   assign dst03 = stage03[60:59];
   assign dst04 = stage04[70:70];
   assign dst05 = stage05[61:60];
   assign dst06 = stage06[51:50];
   assign dst07 = stage07[61:60];
   assign dst08 = stage08[56:55];
   assign dst09 = stage09[70:69];
   assign dst10 = stage10[62:61];
   assign dst11 = stage11[56:55];
   assign dst12 = stage12[57:56];
   assign dst13 = stage13[60:59];
   assign dst14 = stage14[59:58];
   assign dst15 = stage15[57:56];
   assign dst16 = stage16[66:65];
   assign dst17 = stage17[54:53];
   assign dst18 = stage18[57:56];
   assign dst19 = stage19[60:59];
   assign dst20 = stage20[58:57];
   assign dst21 = stage21[57:56];
   assign dst22 = stage22[60:59];
   assign dst23 = stage23[63:62];
   assign dst24 = stage24[62:61];
   assign dst25 = stage25[60:59];
   assign dst26 = stage26[67:66];
   assign dst27 = stage27[70:69];
   assign dst28 = stage28[66:65];
   assign dst29 = stage29[61:60];
   assign dst30 = stage30[66:65];
   assign dst31 = stage31[70:69];
   assign dst32 = stage32[17:16];
   assign dst33 = stage33[14:13];
   assign dst34 = stage34[4:3];
   assign dst35 = stage35[2:2];
   assign dst36 = stage36[0:0];
   gpc1_1 gpc1_1_0(
      {stage00[0]},
      {stage00[32]}
   );
   gpc1_1 gpc1_1_1(
      {stage00[1]},
      {stage00[33]}
   );
   gpc1_1 gpc1_1_2(
      {stage00[2]},
      {stage00[34]}
   );
   gpc1_1 gpc1_1_3(
      {stage00[3]},
      {stage00[35]}
   );
   gpc1_1 gpc1_1_4(
      {stage00[4]},
      {stage00[36]}
   );
   gpc1_1 gpc1_1_5(
      {stage00[5]},
      {stage00[37]}
   );
   gpc1_1 gpc1_1_6(
      {stage00[6]},
      {stage00[38]}
   );
   gpc615_5 gpc615_5_7(
      {stage00[7], stage00[8], stage00[9], stage00[10], stage00[11]},
      {stage01[0]},
      {stage02[0], stage02[1], stage02[2], stage02[3], stage02[4], stage02[5]},
      {stage04[32], stage03[32], stage02[32], stage01[32], stage00[39]}
   );
   gpc615_5 gpc615_5_8(
      {stage00[12], stage00[13], stage00[14], stage00[15], stage00[16]},
      {stage01[1]},
      {stage02[6], stage02[7], stage02[8], stage02[9], stage02[10], stage02[11]},
      {stage04[33], stage03[33], stage02[33], stage01[33], stage00[40]}
   );
   gpc615_5 gpc615_5_9(
      {stage00[17], stage00[18], stage00[19], stage00[20], stage00[21]},
      {stage01[2]},
      {stage02[12], stage02[13], stage02[14], stage02[15], stage02[16], stage02[17]},
      {stage04[34], stage03[34], stage02[34], stage01[34], stage00[41]}
   );
   gpc615_5 gpc615_5_10(
      {stage00[22], stage00[23], stage00[24], stage00[25], stage00[26]},
      {stage01[3]},
      {stage02[18], stage02[19], stage02[20], stage02[21], stage02[22], stage02[23]},
      {stage04[35], stage03[35], stage02[35], stage01[35], stage00[42]}
   );
   gpc615_5 gpc615_5_11(
      {stage00[27], stage00[28], stage00[29], stage00[30], stage00[31]},
      {stage01[4]},
      {stage02[24], stage02[25], stage02[26], stage02[27], stage02[28], stage02[29]},
      {stage04[36], stage03[36], stage02[36], stage01[36], stage00[43]}
   );
   gpc1_1 gpc1_1_12(
      {stage01[5]},
      {stage01[37]}
   );
   gpc1_1 gpc1_1_13(
      {stage01[6]},
      {stage01[38]}
   );
   gpc1_1 gpc1_1_14(
      {stage01[7]},
      {stage01[39]}
   );
   gpc606_5 gpc606_5_15(
      {stage01[8], stage01[9], stage01[10], stage01[11], stage01[12], stage01[13]},
      {stage03[0], stage03[1], stage03[2], stage03[3], stage03[4], stage03[5]},
      {stage05[32], stage04[37], stage03[37], stage02[37], stage01[40]}
   );
   gpc606_5 gpc606_5_16(
      {stage01[14], stage01[15], stage01[16], stage01[17], stage01[18], stage01[19]},
      {stage03[6], stage03[7], stage03[8], stage03[9], stage03[10], stage03[11]},
      {stage05[33], stage04[38], stage03[38], stage02[38], stage01[41]}
   );
   gpc606_5 gpc606_5_17(
      {stage01[20], stage01[21], stage01[22], stage01[23], stage01[24], stage01[25]},
      {stage03[12], stage03[13], stage03[14], stage03[15], stage03[16], stage03[17]},
      {stage05[34], stage04[39], stage03[39], stage02[39], stage01[42]}
   );
   gpc606_5 gpc606_5_18(
      {stage01[26], stage01[27], stage01[28], stage01[29], stage01[30], stage01[31]},
      {stage03[18], stage03[19], stage03[20], stage03[21], stage03[22], stage03[23]},
      {stage05[35], stage04[40], stage03[40], stage02[40], stage01[43]}
   );
   gpc1_1 gpc1_1_19(
      {stage02[30]},
      {stage02[41]}
   );
   gpc1_1 gpc1_1_20(
      {stage02[31]},
      {stage02[42]}
   );
   gpc1_1 gpc1_1_21(
      {stage03[24]},
      {stage03[41]}
   );
   gpc1_1 gpc1_1_22(
      {stage03[25]},
      {stage03[42]}
   );
   gpc1_1 gpc1_1_23(
      {stage03[26]},
      {stage03[43]}
   );
   gpc1_1 gpc1_1_24(
      {stage03[27]},
      {stage03[44]}
   );
   gpc1_1 gpc1_1_25(
      {stage03[28]},
      {stage03[45]}
   );
   gpc1_1 gpc1_1_26(
      {stage03[29]},
      {stage03[46]}
   );
   gpc1_1 gpc1_1_27(
      {stage03[30]},
      {stage03[47]}
   );
   gpc1_1 gpc1_1_28(
      {stage03[31]},
      {stage03[48]}
   );
   gpc1_1 gpc1_1_29(
      {stage04[0]},
      {stage04[41]}
   );
   gpc1_1 gpc1_1_30(
      {stage04[1]},
      {stage04[42]}
   );
   gpc1_1 gpc1_1_31(
      {stage04[2]},
      {stage04[43]}
   );
   gpc1_1 gpc1_1_32(
      {stage04[3]},
      {stage04[44]}
   );
   gpc1_1 gpc1_1_33(
      {stage04[4]},
      {stage04[45]}
   );
   gpc1_1 gpc1_1_34(
      {stage04[5]},
      {stage04[46]}
   );
   gpc1_1 gpc1_1_35(
      {stage04[6]},
      {stage04[47]}
   );
   gpc1_1 gpc1_1_36(
      {stage04[7]},
      {stage04[48]}
   );
   gpc1_1 gpc1_1_37(
      {stage04[8]},
      {stage04[49]}
   );
   gpc606_5 gpc606_5_38(
      {stage04[9], stage04[10], stage04[11], stage04[12], stage04[13], stage04[14]},
      {stage06[0], stage06[1], stage06[2], stage06[3], stage06[4], stage06[5]},
      {stage08[32], stage07[32], stage06[32], stage05[36], stage04[50]}
   );
   gpc606_5 gpc606_5_39(
      {stage04[15], stage04[16], stage04[17], stage04[18], stage04[19], stage04[20]},
      {stage06[6], stage06[7], stage06[8], stage06[9], stage06[10], stage06[11]},
      {stage08[33], stage07[33], stage06[33], stage05[37], stage04[51]}
   );
   gpc606_5 gpc606_5_40(
      {stage04[21], stage04[22], stage04[23], stage04[24], stage04[25], stage04[26]},
      {stage06[12], stage06[13], stage06[14], stage06[15], stage06[16], stage06[17]},
      {stage08[34], stage07[34], stage06[34], stage05[38], stage04[52]}
   );
   gpc1325_5 gpc1325_5_41(
      {stage04[27], stage04[28], stage04[29], stage04[30], stage04[31]},
      {stage05[0], stage05[1]},
      {stage06[18], stage06[19], stage06[20]},
      {stage07[0]},
      {stage08[35], stage07[35], stage06[35], stage05[39], stage04[53]}
   );
   gpc1_1 gpc1_1_42(
      {stage05[2]},
      {stage05[40]}
   );
   gpc1_1 gpc1_1_43(
      {stage05[3]},
      {stage05[41]}
   );
   gpc1_1 gpc1_1_44(
      {stage05[4]},
      {stage05[42]}
   );
   gpc1_1 gpc1_1_45(
      {stage05[5]},
      {stage05[43]}
   );
   gpc1_1 gpc1_1_46(
      {stage05[6]},
      {stage05[44]}
   );
   gpc1_1 gpc1_1_47(
      {stage05[7]},
      {stage05[45]}
   );
   gpc606_5 gpc606_5_48(
      {stage05[8], stage05[9], stage05[10], stage05[11], stage05[12], stage05[13]},
      {stage07[1], stage07[2], stage07[3], stage07[4], stage07[5], stage07[6]},
      {stage09[32], stage08[36], stage07[36], stage06[36], stage05[46]}
   );
   gpc606_5 gpc606_5_49(
      {stage05[14], stage05[15], stage05[16], stage05[17], stage05[18], stage05[19]},
      {stage07[7], stage07[8], stage07[9], stage07[10], stage07[11], stage07[12]},
      {stage09[33], stage08[37], stage07[37], stage06[37], stage05[47]}
   );
   gpc606_5 gpc606_5_50(
      {stage05[20], stage05[21], stage05[22], stage05[23], stage05[24], stage05[25]},
      {stage07[13], stage07[14], stage07[15], stage07[16], stage07[17], stage07[18]},
      {stage09[34], stage08[38], stage07[38], stage06[38], stage05[48]}
   );
   gpc606_5 gpc606_5_51(
      {stage05[26], stage05[27], stage05[28], stage05[29], stage05[30], stage05[31]},
      {stage07[19], stage07[20], stage07[21], stage07[22], stage07[23], stage07[24]},
      {stage09[35], stage08[39], stage07[39], stage06[39], stage05[49]}
   );
   gpc606_5 gpc606_5_52(
      {stage06[21], stage06[22], stage06[23], stage06[24], stage06[25], stage06[26]},
      {stage08[0], stage08[1], stage08[2], stage08[3], stage08[4], stage08[5]},
      {stage10[32], stage09[36], stage08[40], stage07[40], stage06[40]}
   );
   gpc615_5 gpc615_5_53(
      {stage06[27], stage06[28], stage06[29], stage06[30], stage06[31]},
      {stage07[25]},
      {stage08[6], stage08[7], stage08[8], stage08[9], stage08[10], stage08[11]},
      {stage10[33], stage09[37], stage08[41], stage07[41], stage06[41]}
   );
   gpc1_1 gpc1_1_54(
      {stage07[26]},
      {stage07[42]}
   );
   gpc1_1 gpc1_1_55(
      {stage07[27]},
      {stage07[43]}
   );
   gpc1_1 gpc1_1_56(
      {stage07[28]},
      {stage07[44]}
   );
   gpc623_5 gpc623_5_57(
      {stage07[29], stage07[30], stage07[31]},
      {stage08[12], stage08[13]},
      {stage09[0], stage09[1], stage09[2], stage09[3], stage09[4], stage09[5]},
      {stage11[32], stage10[34], stage09[38], stage08[42], stage07[45]}
   );
   gpc606_5 gpc606_5_58(
      {stage08[14], stage08[15], stage08[16], stage08[17], stage08[18], stage08[19]},
      {stage10[0], stage10[1], stage10[2], stage10[3], stage10[4], stage10[5]},
      {stage12[32], stage11[33], stage10[35], stage09[39], stage08[43]}
   );
   gpc606_5 gpc606_5_59(
      {stage08[20], stage08[21], stage08[22], stage08[23], stage08[24], stage08[25]},
      {stage10[6], stage10[7], stage10[8], stage10[9], stage10[10], stage10[11]},
      {stage12[33], stage11[34], stage10[36], stage09[40], stage08[44]}
   );
   gpc606_5 gpc606_5_60(
      {stage08[26], stage08[27], stage08[28], stage08[29], stage08[30], stage08[31]},
      {stage10[12], stage10[13], stage10[14], stage10[15], stage10[16], stage10[17]},
      {stage12[34], stage11[35], stage10[37], stage09[41], stage08[45]}
   );
   gpc1_1 gpc1_1_61(
      {stage09[6]},
      {stage09[42]}
   );
   gpc1_1 gpc1_1_62(
      {stage09[7]},
      {stage09[43]}
   );
   gpc1_1 gpc1_1_63(
      {stage09[8]},
      {stage09[44]}
   );
   gpc1_1 gpc1_1_64(
      {stage09[9]},
      {stage09[45]}
   );
   gpc1_1 gpc1_1_65(
      {stage09[10]},
      {stage09[46]}
   );
   gpc1_1 gpc1_1_66(
      {stage09[11]},
      {stage09[47]}
   );
   gpc1_1 gpc1_1_67(
      {stage09[12]},
      {stage09[48]}
   );
   gpc1_1 gpc1_1_68(
      {stage09[13]},
      {stage09[49]}
   );
   gpc606_5 gpc606_5_69(
      {stage09[14], stage09[15], stage09[16], stage09[17], stage09[18], stage09[19]},
      {stage11[0], stage11[1], stage11[2], stage11[3], stage11[4], stage11[5]},
      {stage13[32], stage12[35], stage11[36], stage10[38], stage09[50]}
   );
   gpc606_5 gpc606_5_70(
      {stage09[20], stage09[21], stage09[22], stage09[23], stage09[24], stage09[25]},
      {stage11[6], stage11[7], stage11[8], stage11[9], stage11[10], stage11[11]},
      {stage13[33], stage12[36], stage11[37], stage10[39], stage09[51]}
   );
   gpc606_5 gpc606_5_71(
      {stage09[26], stage09[27], stage09[28], stage09[29], stage09[30], stage09[31]},
      {stage11[12], stage11[13], stage11[14], stage11[15], stage11[16], stage11[17]},
      {stage13[34], stage12[37], stage11[38], stage10[40], stage09[52]}
   );
   gpc1_1 gpc1_1_72(
      {stage10[18]},
      {stage10[41]}
   );
   gpc1_1 gpc1_1_73(
      {stage10[19]},
      {stage10[42]}
   );
   gpc1_1 gpc1_1_74(
      {stage10[20]},
      {stage10[43]}
   );
   gpc1_1 gpc1_1_75(
      {stage10[21]},
      {stage10[44]}
   );
   gpc615_5 gpc615_5_76(
      {stage10[22], stage10[23], stage10[24], stage10[25], stage10[26]},
      {stage11[18]},
      {stage12[0], stage12[1], stage12[2], stage12[3], stage12[4], stage12[5]},
      {stage14[32], stage13[35], stage12[38], stage11[39], stage10[45]}
   );
   gpc615_5 gpc615_5_77(
      {stage10[27], stage10[28], stage10[29], stage10[30], stage10[31]},
      {stage11[19]},
      {stage12[6], stage12[7], stage12[8], stage12[9], stage12[10], stage12[11]},
      {stage14[33], stage13[36], stage12[39], stage11[40], stage10[46]}
   );
   gpc1_1 gpc1_1_78(
      {stage11[20]},
      {stage11[41]}
   );
   gpc1_1 gpc1_1_79(
      {stage11[21]},
      {stage11[42]}
   );
   gpc615_5 gpc615_5_80(
      {stage11[22], stage11[23], stage11[24], stage11[25], stage11[26]},
      {stage12[12]},
      {stage13[0], stage13[1], stage13[2], stage13[3], stage13[4], stage13[5]},
      {stage15[32], stage14[34], stage13[37], stage12[40], stage11[43]}
   );
   gpc615_5 gpc615_5_81(
      {stage11[27], stage11[28], stage11[29], stage11[30], stage11[31]},
      {stage12[13]},
      {stage13[6], stage13[7], stage13[8], stage13[9], stage13[10], stage13[11]},
      {stage15[33], stage14[35], stage13[38], stage12[41], stage11[44]}
   );
   gpc1_1 gpc1_1_82(
      {stage12[14]},
      {stage12[42]}
   );
   gpc606_5 gpc606_5_83(
      {stage12[15], stage12[16], stage12[17], stage12[18], stage12[19], stage12[20]},
      {stage14[0], stage14[1], stage14[2], stage14[3], stage14[4], stage14[5]},
      {stage16[32], stage15[34], stage14[36], stage13[39], stage12[43]}
   );
   gpc606_5 gpc606_5_84(
      {stage12[21], stage12[22], stage12[23], stage12[24], stage12[25], stage12[26]},
      {stage14[6], stage14[7], stage14[8], stage14[9], stage14[10], stage14[11]},
      {stage16[33], stage15[35], stage14[37], stage13[40], stage12[44]}
   );
   gpc615_5 gpc615_5_85(
      {stage12[27], stage12[28], stage12[29], stage12[30], stage12[31]},
      {stage13[12]},
      {stage14[12], stage14[13], stage14[14], stage14[15], stage14[16], stage14[17]},
      {stage16[34], stage15[36], stage14[38], stage13[41], stage12[45]}
   );
   gpc1_1 gpc1_1_86(
      {stage13[13]},
      {stage13[42]}
   );
   gpc1_1 gpc1_1_87(
      {stage13[14]},
      {stage13[43]}
   );
   gpc1_1 gpc1_1_88(
      {stage13[15]},
      {stage13[44]}
   );
   gpc606_5 gpc606_5_89(
      {stage13[16], stage13[17], stage13[18], stage13[19], stage13[20], stage13[21]},
      {stage15[0], stage15[1], stage15[2], stage15[3], stage15[4], stage15[5]},
      {stage17[32], stage16[35], stage15[37], stage14[39], stage13[45]}
   );
   gpc615_5 gpc615_5_90(
      {stage13[22], stage13[23], stage13[24], stage13[25], stage13[26]},
      {stage14[18]},
      {stage15[6], stage15[7], stage15[8], stage15[9], stage15[10], stage15[11]},
      {stage17[33], stage16[36], stage15[38], stage14[40], stage13[46]}
   );
   gpc615_5 gpc615_5_91(
      {stage13[27], stage13[28], stage13[29], stage13[30], stage13[31]},
      {stage14[19]},
      {stage15[12], stage15[13], stage15[14], stage15[15], stage15[16], stage15[17]},
      {stage17[34], stage16[37], stage15[39], stage14[41], stage13[47]}
   );
   gpc1_1 gpc1_1_92(
      {stage14[20]},
      {stage14[42]}
   );
   gpc1_1 gpc1_1_93(
      {stage14[21]},
      {stage14[43]}
   );
   gpc1_1 gpc1_1_94(
      {stage14[22]},
      {stage14[44]}
   );
   gpc1_1 gpc1_1_95(
      {stage14[23]},
      {stage14[45]}
   );
   gpc1_1 gpc1_1_96(
      {stage14[24]},
      {stage14[46]}
   );
   gpc1_1 gpc1_1_97(
      {stage14[25]},
      {stage14[47]}
   );
   gpc1_1 gpc1_1_98(
      {stage14[26]},
      {stage14[48]}
   );
   gpc615_5 gpc615_5_99(
      {stage14[27], stage14[28], stage14[29], stage14[30], stage14[31]},
      {stage15[18]},
      {stage16[0], stage16[1], stage16[2], stage16[3], stage16[4], stage16[5]},
      {stage18[32], stage17[35], stage16[38], stage15[40], stage14[49]}
   );
   gpc615_5 gpc615_5_100(
      {stage15[19], stage15[20], stage15[21], stage15[22], stage15[23]},
      {stage16[6]},
      {stage17[0], stage17[1], stage17[2], stage17[3], stage17[4], stage17[5]},
      {stage19[32], stage18[33], stage17[36], stage16[39], stage15[41]}
   );
   gpc615_5 gpc615_5_101(
      {stage15[24], stage15[25], stage15[26], stage15[27], stage15[28]},
      {stage16[7]},
      {stage17[6], stage17[7], stage17[8], stage17[9], stage17[10], stage17[11]},
      {stage19[33], stage18[34], stage17[37], stage16[40], stage15[42]}
   );
   gpc1325_5 gpc1325_5_102(
      {stage15[29], stage15[30], stage15[31], 1'h0, 1'h0},
      {stage16[8], stage16[9]},
      {stage17[12], stage17[13], stage17[14]},
      {stage18[0]},
      {stage19[34], stage18[35], stage17[38], stage16[41], stage15[43]}
   );
   gpc1_1 gpc1_1_103(
      {stage16[10]},
      {stage16[42]}
   );
   gpc1_1 gpc1_1_104(
      {stage16[11]},
      {stage16[43]}
   );
   gpc1_1 gpc1_1_105(
      {stage16[12]},
      {stage16[44]}
   );
   gpc1_1 gpc1_1_106(
      {stage16[13]},
      {stage16[45]}
   );
   gpc1_1 gpc1_1_107(
      {stage16[14]},
      {stage16[46]}
   );
   gpc606_5 gpc606_5_108(
      {stage16[15], stage16[16], stage16[17], stage16[18], stage16[19], stage16[20]},
      {stage18[1], stage18[2], stage18[3], stage18[4], stage18[5], stage18[6]},
      {stage20[32], stage19[35], stage18[36], stage17[39], stage16[47]}
   );
   gpc606_5 gpc606_5_109(
      {stage16[21], stage16[22], stage16[23], stage16[24], stage16[25], stage16[26]},
      {stage18[7], stage18[8], stage18[9], stage18[10], stage18[11], stage18[12]},
      {stage20[33], stage19[36], stage18[37], stage17[40], stage16[48]}
   );
   gpc615_5 gpc615_5_110(
      {stage16[27], stage16[28], stage16[29], stage16[30], stage16[31]},
      {stage17[15]},
      {stage18[13], stage18[14], stage18[15], stage18[16], stage18[17], stage18[18]},
      {stage20[34], stage19[37], stage18[38], stage17[41], stage16[49]}
   );
   gpc606_5 gpc606_5_111(
      {stage17[16], stage17[17], stage17[18], stage17[19], stage17[20], stage17[21]},
      {stage19[0], stage19[1], stage19[2], stage19[3], stage19[4], stage19[5]},
      {stage21[32], stage20[35], stage19[38], stage18[39], stage17[42]}
   );
   gpc615_5 gpc615_5_112(
      {stage17[22], stage17[23], stage17[24], stage17[25], stage17[26]},
      {stage18[19]},
      {stage19[6], stage19[7], stage19[8], stage19[9], stage19[10], stage19[11]},
      {stage21[33], stage20[36], stage19[39], stage18[40], stage17[43]}
   );
   gpc2135_5 gpc2135_5_113(
      {stage17[27], stage17[28], stage17[29], stage17[30], stage17[31]},
      {stage18[20], stage18[21], stage18[22]},
      {stage19[12]},
      {stage20[0], stage20[1]},
      {stage21[34], stage20[37], stage19[40], stage18[41], stage17[44]}
   );
   gpc615_5 gpc615_5_114(
      {stage18[23], stage18[24], stage18[25], stage18[26], stage18[27]},
      {stage19[13]},
      {stage20[2], stage20[3], stage20[4], stage20[5], stage20[6], stage20[7]},
      {stage22[32], stage21[35], stage20[38], stage19[41], stage18[42]}
   );
   gpc615_5 gpc615_5_115(
      {stage18[28], stage18[29], stage18[30], stage18[31], 1'h0},
      {stage19[14]},
      {stage20[8], stage20[9], stage20[10], stage20[11], stage20[12], stage20[13]},
      {stage22[33], stage21[36], stage20[39], stage19[42], stage18[43]}
   );
   gpc1_1 gpc1_1_116(
      {stage19[15]},
      {stage19[43]}
   );
   gpc606_5 gpc606_5_117(
      {stage19[16], stage19[17], stage19[18], stage19[19], stage19[20], stage19[21]},
      {stage21[0], stage21[1], stage21[2], stage21[3], stage21[4], stage21[5]},
      {stage23[32], stage22[34], stage21[37], stage20[40], stage19[44]}
   );
   gpc615_5 gpc615_5_118(
      {stage19[22], stage19[23], stage19[24], stage19[25], stage19[26]},
      {stage20[14]},
      {stage21[6], stage21[7], stage21[8], stage21[9], stage21[10], stage21[11]},
      {stage23[33], stage22[35], stage21[38], stage20[41], stage19[45]}
   );
   gpc615_5 gpc615_5_119(
      {stage19[27], stage19[28], stage19[29], stage19[30], stage19[31]},
      {stage20[15]},
      {stage21[12], stage21[13], stage21[14], stage21[15], stage21[16], stage21[17]},
      {stage23[34], stage22[36], stage21[39], stage20[42], stage19[46]}
   );
   gpc1_1 gpc1_1_120(
      {stage20[16]},
      {stage20[43]}
   );
   gpc1_1 gpc1_1_121(
      {stage20[17]},
      {stage20[44]}
   );
   gpc1_1 gpc1_1_122(
      {stage20[18]},
      {stage20[45]}
   );
   gpc1_1 gpc1_1_123(
      {stage20[19]},
      {stage20[46]}
   );
   gpc606_5 gpc606_5_124(
      {stage20[20], stage20[21], stage20[22], stage20[23], stage20[24], stage20[25]},
      {stage22[0], stage22[1], stage22[2], stage22[3], stage22[4], stage22[5]},
      {stage24[32], stage23[35], stage22[37], stage21[40], stage20[47]}
   );
   gpc606_5 gpc606_5_125(
      {stage20[26], stage20[27], stage20[28], stage20[29], stage20[30], stage20[31]},
      {stage22[6], stage22[7], stage22[8], stage22[9], stage22[10], stage22[11]},
      {stage24[33], stage23[36], stage22[38], stage21[41], stage20[48]}
   );
   gpc1_1 gpc1_1_126(
      {stage21[18]},
      {stage21[42]}
   );
   gpc1_1 gpc1_1_127(
      {stage21[19]},
      {stage21[43]}
   );
   gpc1_1 gpc1_1_128(
      {stage21[20]},
      {stage21[44]}
   );
   gpc1_1 gpc1_1_129(
      {stage21[21]},
      {stage21[45]}
   );
   gpc615_5 gpc615_5_130(
      {stage21[22], stage21[23], stage21[24], stage21[25], stage21[26]},
      {stage22[12]},
      {stage23[0], stage23[1], stage23[2], stage23[3], stage23[4], stage23[5]},
      {stage25[32], stage24[34], stage23[37], stage22[39], stage21[46]}
   );
   gpc615_5 gpc615_5_131(
      {stage21[27], stage21[28], stage21[29], stage21[30], stage21[31]},
      {stage22[13]},
      {stage23[6], stage23[7], stage23[8], stage23[9], stage23[10], stage23[11]},
      {stage25[33], stage24[35], stage23[38], stage22[40], stage21[47]}
   );
   gpc1_1 gpc1_1_132(
      {stage22[14]},
      {stage22[41]}
   );
   gpc1_1 gpc1_1_133(
      {stage22[15]},
      {stage22[42]}
   );
   gpc1_1 gpc1_1_134(
      {stage22[16]},
      {stage22[43]}
   );
   gpc615_5 gpc615_5_135(
      {stage22[17], stage22[18], stage22[19], stage22[20], stage22[21]},
      {stage23[12]},
      {stage24[0], stage24[1], stage24[2], stage24[3], stage24[4], stage24[5]},
      {stage26[32], stage25[34], stage24[36], stage23[39], stage22[44]}
   );
   gpc615_5 gpc615_5_136(
      {stage22[22], stage22[23], stage22[24], stage22[25], stage22[26]},
      {stage23[13]},
      {stage24[6], stage24[7], stage24[8], stage24[9], stage24[10], stage24[11]},
      {stage26[33], stage25[35], stage24[37], stage23[40], stage22[45]}
   );
   gpc2135_5 gpc2135_5_137(
      {stage22[27], stage22[28], stage22[29], stage22[30], stage22[31]},
      {stage23[14], stage23[15], stage23[16]},
      {stage24[12]},
      {stage25[0], stage25[1]},
      {stage26[34], stage25[36], stage24[38], stage23[41], stage22[46]}
   );
   gpc1_1 gpc1_1_138(
      {stage23[17]},
      {stage23[42]}
   );
   gpc1_1 gpc1_1_139(
      {stage23[18]},
      {stage23[43]}
   );
   gpc1_1 gpc1_1_140(
      {stage23[19]},
      {stage23[44]}
   );
   gpc1_1 gpc1_1_141(
      {stage23[20]},
      {stage23[45]}
   );
   gpc1_1 gpc1_1_142(
      {stage23[21]},
      {stage23[46]}
   );
   gpc615_5 gpc615_5_143(
      {stage23[22], stage23[23], stage23[24], stage23[25], stage23[26]},
      {stage24[13]},
      {stage25[2], stage25[3], stage25[4], stage25[5], stage25[6], stage25[7]},
      {stage27[32], stage26[35], stage25[37], stage24[39], stage23[47]}
   );
   gpc615_5 gpc615_5_144(
      {stage23[27], stage23[28], stage23[29], stage23[30], stage23[31]},
      {stage24[14]},
      {stage25[8], stage25[9], stage25[10], stage25[11], stage25[12], stage25[13]},
      {stage27[33], stage26[36], stage25[38], stage24[40], stage23[48]}
   );
   gpc1_1 gpc1_1_145(
      {stage24[15]},
      {stage24[41]}
   );
   gpc1_1 gpc1_1_146(
      {stage24[16]},
      {stage24[42]}
   );
   gpc1_1 gpc1_1_147(
      {stage24[17]},
      {stage24[43]}
   );
   gpc1_1 gpc1_1_148(
      {stage24[18]},
      {stage24[44]}
   );
   gpc1_1 gpc1_1_149(
      {stage24[19]},
      {stage24[45]}
   );
   gpc1_1 gpc1_1_150(
      {stage24[20]},
      {stage24[46]}
   );
   gpc1_1 gpc1_1_151(
      {stage24[21]},
      {stage24[47]}
   );
   gpc615_5 gpc615_5_152(
      {stage24[22], stage24[23], stage24[24], stage24[25], stage24[26]},
      {stage25[14]},
      {stage26[0], stage26[1], stage26[2], stage26[3], stage26[4], stage26[5]},
      {stage28[32], stage27[34], stage26[37], stage25[39], stage24[48]}
   );
   gpc615_5 gpc615_5_153(
      {stage24[27], stage24[28], stage24[29], stage24[30], stage24[31]},
      {stage25[15]},
      {stage26[6], stage26[7], stage26[8], stage26[9], stage26[10], stage26[11]},
      {stage28[33], stage27[35], stage26[38], stage25[40], stage24[49]}
   );
   gpc615_5 gpc615_5_154(
      {stage25[16], stage25[17], stage25[18], stage25[19], stage25[20]},
      {stage26[12]},
      {stage27[0], stage27[1], stage27[2], stage27[3], stage27[4], stage27[5]},
      {stage29[32], stage28[34], stage27[36], stage26[39], stage25[41]}
   );
   gpc615_5 gpc615_5_155(
      {stage25[21], stage25[22], stage25[23], stage25[24], stage25[25]},
      {stage26[13]},
      {stage27[6], stage27[7], stage27[8], stage27[9], stage27[10], stage27[11]},
      {stage29[33], stage28[35], stage27[37], stage26[40], stage25[42]}
   );
   gpc1343_5 gpc1343_5_156(
      {stage25[26], stage25[27], stage25[28]},
      {stage26[14], stage26[15], stage26[16], stage26[17]},
      {stage27[12], stage27[13], stage27[14]},
      {stage28[0]},
      {stage29[34], stage28[36], stage27[38], stage26[41], stage25[43]}
   );
   gpc1343_5 gpc1343_5_157(
      {stage25[29], stage25[30], stage25[31]},
      {stage26[18], stage26[19], stage26[20], stage26[21]},
      {stage27[15], stage27[16], stage27[17]},
      {stage28[1]},
      {stage29[35], stage28[37], stage27[39], stage26[42], stage25[44]}
   );
   gpc1_1 gpc1_1_158(
      {stage26[22]},
      {stage26[43]}
   );
   gpc1_1 gpc1_1_159(
      {stage26[23]},
      {stage26[44]}
   );
   gpc1_1 gpc1_1_160(
      {stage26[24]},
      {stage26[45]}
   );
   gpc1_1 gpc1_1_161(
      {stage26[25]},
      {stage26[46]}
   );
   gpc1_1 gpc1_1_162(
      {stage26[26]},
      {stage26[47]}
   );
   gpc1_1 gpc1_1_163(
      {stage26[27]},
      {stage26[48]}
   );
   gpc1_1 gpc1_1_164(
      {stage26[28]},
      {stage26[49]}
   );
   gpc1_1 gpc1_1_165(
      {stage26[29]},
      {stage26[50]}
   );
   gpc1_1 gpc1_1_166(
      {stage26[30]},
      {stage26[51]}
   );
   gpc1_1 gpc1_1_167(
      {stage26[31]},
      {stage26[52]}
   );
   gpc1_1 gpc1_1_168(
      {stage27[18]},
      {stage27[40]}
   );
   gpc1_1 gpc1_1_169(
      {stage27[19]},
      {stage27[41]}
   );
   gpc1_1 gpc1_1_170(
      {stage27[20]},
      {stage27[42]}
   );
   gpc1_1 gpc1_1_171(
      {stage27[21]},
      {stage27[43]}
   );
   gpc1_1 gpc1_1_172(
      {stage27[22]},
      {stage27[44]}
   );
   gpc1_1 gpc1_1_173(
      {stage27[23]},
      {stage27[45]}
   );
   gpc1_1 gpc1_1_174(
      {stage27[24]},
      {stage27[46]}
   );
   gpc1_1 gpc1_1_175(
      {stage27[25]},
      {stage27[47]}
   );
   gpc1_1 gpc1_1_176(
      {stage27[26]},
      {stage27[48]}
   );
   gpc1325_5 gpc1325_5_177(
      {stage27[27], stage27[28], stage27[29], stage27[30], stage27[31]},
      {stage28[2], stage28[3]},
      {stage29[0], stage29[1], stage29[2]},
      {stage30[0]},
      {stage31[32], stage30[32], stage29[36], stage28[38], stage27[49]}
   );
   gpc1_1 gpc1_1_178(
      {stage28[4]},
      {stage28[39]}
   );
   gpc1_1 gpc1_1_179(
      {stage28[5]},
      {stage28[40]}
   );
   gpc1_1 gpc1_1_180(
      {stage28[6]},
      {stage28[41]}
   );
   gpc1_1 gpc1_1_181(
      {stage28[7]},
      {stage28[42]}
   );
   gpc1_1 gpc1_1_182(
      {stage28[8]},
      {stage28[43]}
   );
   gpc1_1 gpc1_1_183(
      {stage28[9]},
      {stage28[44]}
   );
   gpc1_1 gpc1_1_184(
      {stage28[10]},
      {stage28[45]}
   );
   gpc1_1 gpc1_1_185(
      {stage28[11]},
      {stage28[46]}
   );
   gpc1_1 gpc1_1_186(
      {stage28[12]},
      {stage28[47]}
   );
   gpc1_1 gpc1_1_187(
      {stage28[13]},
      {stage28[48]}
   );
   gpc1_1 gpc1_1_188(
      {stage28[14]},
      {stage28[49]}
   );
   gpc1_1 gpc1_1_189(
      {stage28[15]},
      {stage28[50]}
   );
   gpc1_1 gpc1_1_190(
      {stage28[16]},
      {stage28[51]}
   );
   gpc615_5 gpc615_5_191(
      {stage28[17], stage28[18], stage28[19], stage28[20], stage28[21]},
      {stage29[3]},
      {stage30[1], stage30[2], stage30[3], stage30[4], stage30[5], stage30[6]},
      {stage32[0], stage31[33], stage30[33], stage29[37], stage28[52]}
   );
   gpc615_5 gpc615_5_192(
      {stage28[22], stage28[23], stage28[24], stage28[25], stage28[26]},
      {stage29[4]},
      {stage30[7], stage30[8], stage30[9], stage30[10], stage30[11], stage30[12]},
      {stage32[1], stage31[34], stage30[34], stage29[38], stage28[53]}
   );
   gpc615_5 gpc615_5_193(
      {stage28[27], stage28[28], stage28[29], stage28[30], stage28[31]},
      {stage29[5]},
      {stage30[13], stage30[14], stage30[15], stage30[16], stage30[17], stage30[18]},
      {stage32[2], stage31[35], stage30[35], stage29[39], stage28[54]}
   );
   gpc1_1 gpc1_1_194(
      {stage29[6]},
      {stage29[40]}
   );
   gpc1_1 gpc1_1_195(
      {stage29[7]},
      {stage29[41]}
   );
   gpc606_5 gpc606_5_196(
      {stage29[8], stage29[9], stage29[10], stage29[11], stage29[12], stage29[13]},
      {stage31[0], stage31[1], stage31[2], stage31[3], stage31[4], stage31[5]},
      {stage33[0], stage32[3], stage31[36], stage30[36], stage29[42]}
   );
   gpc606_5 gpc606_5_197(
      {stage29[14], stage29[15], stage29[16], stage29[17], stage29[18], stage29[19]},
      {stage31[6], stage31[7], stage31[8], stage31[9], stage31[10], stage31[11]},
      {stage33[1], stage32[4], stage31[37], stage30[37], stage29[43]}
   );
   gpc606_5 gpc606_5_198(
      {stage29[20], stage29[21], stage29[22], stage29[23], stage29[24], stage29[25]},
      {stage31[12], stage31[13], stage31[14], stage31[15], stage31[16], stage31[17]},
      {stage33[2], stage32[5], stage31[38], stage30[38], stage29[44]}
   );
   gpc606_5 gpc606_5_199(
      {stage29[26], stage29[27], stage29[28], stage29[29], stage29[30], stage29[31]},
      {stage31[18], stage31[19], stage31[20], stage31[21], stage31[22], stage31[23]},
      {stage33[3], stage32[6], stage31[39], stage30[39], stage29[45]}
   );
   gpc1_1 gpc1_1_200(
      {stage30[19]},
      {stage30[40]}
   );
   gpc1_1 gpc1_1_201(
      {stage30[20]},
      {stage30[41]}
   );
   gpc1_1 gpc1_1_202(
      {stage30[21]},
      {stage30[42]}
   );
   gpc1_1 gpc1_1_203(
      {stage30[22]},
      {stage30[43]}
   );
   gpc1_1 gpc1_1_204(
      {stage30[23]},
      {stage30[44]}
   );
   gpc1_1 gpc1_1_205(
      {stage30[24]},
      {stage30[45]}
   );
   gpc1_1 gpc1_1_206(
      {stage30[25]},
      {stage30[46]}
   );
   gpc1_1 gpc1_1_207(
      {stage30[26]},
      {stage30[47]}
   );
   gpc1_1 gpc1_1_208(
      {stage30[27]},
      {stage30[48]}
   );
   gpc1_1 gpc1_1_209(
      {stage30[28]},
      {stage30[49]}
   );
   gpc1_1 gpc1_1_210(
      {stage30[29]},
      {stage30[50]}
   );
   gpc1_1 gpc1_1_211(
      {stage30[30]},
      {stage30[51]}
   );
   gpc1_1 gpc1_1_212(
      {stage30[31]},
      {stage30[52]}
   );
   gpc1_1 gpc1_1_213(
      {stage31[24]},
      {stage31[40]}
   );
   gpc1_1 gpc1_1_214(
      {stage31[25]},
      {stage31[41]}
   );
   gpc1_1 gpc1_1_215(
      {stage31[26]},
      {stage31[42]}
   );
   gpc1_1 gpc1_1_216(
      {stage31[27]},
      {stage31[43]}
   );
   gpc1_1 gpc1_1_217(
      {stage31[28]},
      {stage31[44]}
   );
   gpc1_1 gpc1_1_218(
      {stage31[29]},
      {stage31[45]}
   );
   gpc1_1 gpc1_1_219(
      {stage31[30]},
      {stage31[46]}
   );
   gpc1_1 gpc1_1_220(
      {stage31[31]},
      {stage31[47]}
   );
   gpc1_1 gpc1_1_221(
      {stage00[32]},
      {stage00[44]}
   );
   gpc1_1 gpc1_1_222(
      {stage00[33]},
      {stage00[45]}
   );
   gpc615_5 gpc615_5_223(
      {stage00[34], stage00[35], stage00[36], stage00[37], stage00[38]},
      {stage01[32]},
      {stage02[32], stage02[33], stage02[34], stage02[35], stage02[36], stage02[37]},
      {stage04[54], stage03[49], stage02[43], stage01[44], stage00[46]}
   );
   gpc2135_5 gpc2135_5_224(
      {stage00[39], stage00[40], stage00[41], stage00[42], stage00[43]},
      {stage01[33], stage01[34], stage01[35]},
      {stage02[38]},
      {stage03[32], stage03[33]},
      {stage04[55], stage03[50], stage02[44], stage01[45], stage00[47]}
   );
   gpc606_5 gpc606_5_225(
      {stage01[36], stage01[37], stage01[38], stage01[39], stage01[40], stage01[41]},
      {stage03[34], stage03[35], stage03[36], stage03[37], stage03[38], stage03[39]},
      {stage05[50], stage04[56], stage03[51], stage02[45], stage01[46]}
   );
   gpc606_5 gpc606_5_226(
      {stage01[42], stage01[43], 1'h0, 1'h0, 1'h0, 1'h0},
      {stage03[40], stage03[41], stage03[42], stage03[43], stage03[44], stage03[45]},
      {stage05[51], stage04[57], stage03[52], stage02[46], stage01[47]}
   );
   gpc1_1 gpc1_1_227(
      {stage02[39]},
      {stage02[47]}
   );
   gpc1_1 gpc1_1_228(
      {stage02[40]},
      {stage02[48]}
   );
   gpc1_1 gpc1_1_229(
      {stage02[41]},
      {stage02[49]}
   );
   gpc1_1 gpc1_1_230(
      {stage02[42]},
      {stage02[50]}
   );
   gpc1_1 gpc1_1_231(
      {stage03[46]},
      {stage03[53]}
   );
   gpc1_1 gpc1_1_232(
      {stage03[47]},
      {stage03[54]}
   );
   gpc1_1 gpc1_1_233(
      {stage03[48]},
      {stage03[55]}
   );
   gpc1_1 gpc1_1_234(
      {stage04[32]},
      {stage04[58]}
   );
   gpc1_1 gpc1_1_235(
      {stage04[33]},
      {stage04[59]}
   );
   gpc135_4 gpc135_4_236(
      {stage04[34], stage04[35], stage04[36], stage04[37], stage04[38]},
      {stage05[32], stage05[33], stage05[34]},
      {stage06[32]},
      {stage07[46], stage06[42], stage05[52], stage04[60]}
   );
   gpc135_4 gpc135_4_237(
      {stage04[39], stage04[40], stage04[41], stage04[42], stage04[43]},
      {stage05[35], stage05[36], stage05[37]},
      {stage06[33]},
      {stage07[47], stage06[43], stage05[53], stage04[61]}
   );
   gpc135_4 gpc135_4_238(
      {stage04[44], stage04[45], stage04[46], stage04[47], stage04[48]},
      {stage05[38], stage05[39], stage05[40]},
      {stage06[34]},
      {stage07[48], stage06[44], stage05[54], stage04[62]}
   );
   gpc135_4 gpc135_4_239(
      {stage04[49], stage04[50], stage04[51], stage04[52], stage04[53]},
      {stage05[41], stage05[42], stage05[43]},
      {stage06[35]},
      {stage07[49], stage06[45], stage05[55], stage04[63]}
   );
   gpc606_5 gpc606_5_240(
      {stage05[44], stage05[45], stage05[46], stage05[47], stage05[48], stage05[49]},
      {stage07[32], stage07[33], stage07[34], stage07[35], stage07[36], stage07[37]},
      {stage09[53], stage08[46], stage07[50], stage06[46], stage05[56]}
   );
   gpc606_5 gpc606_5_241(
      {stage06[36], stage06[37], stage06[38], stage06[39], stage06[40], stage06[41]},
      {stage08[32], stage08[33], stage08[34], stage08[35], stage08[36], stage08[37]},
      {stage10[47], stage09[54], stage08[47], stage07[51], stage06[47]}
   );
   gpc1_1 gpc1_1_242(
      {stage07[38]},
      {stage07[52]}
   );
   gpc1_1 gpc1_1_243(
      {stage07[39]},
      {stage07[53]}
   );
   gpc1_1 gpc1_1_244(
      {stage07[40]},
      {stage07[54]}
   );
   gpc615_5 gpc615_5_245(
      {stage07[41], stage07[42], stage07[43], stage07[44], stage07[45]},
      {stage08[38]},
      {stage09[32], stage09[33], stage09[34], stage09[35], stage09[36], stage09[37]},
      {stage11[45], stage10[48], stage09[55], stage08[48], stage07[55]}
   );
   gpc1_1 gpc1_1_246(
      {stage08[39]},
      {stage08[49]}
   );
   gpc1_1 gpc1_1_247(
      {stage08[40]},
      {stage08[50]}
   );
   gpc615_5 gpc615_5_248(
      {stage08[41], stage08[42], stage08[43], stage08[44], stage08[45]},
      {stage09[38]},
      {stage10[32], stage10[33], stage10[34], stage10[35], stage10[36], stage10[37]},
      {stage12[46], stage11[46], stage10[49], stage09[56], stage08[51]}
   );
   gpc1_1 gpc1_1_249(
      {stage09[39]},
      {stage09[57]}
   );
   gpc1_1 gpc1_1_250(
      {stage09[40]},
      {stage09[58]}
   );
   gpc1_1 gpc1_1_251(
      {stage09[41]},
      {stage09[59]}
   );
   gpc1_1 gpc1_1_252(
      {stage09[42]},
      {stage09[60]}
   );
   gpc1_1 gpc1_1_253(
      {stage09[43]},
      {stage09[61]}
   );
   gpc1_1 gpc1_1_254(
      {stage09[44]},
      {stage09[62]}
   );
   gpc1_1 gpc1_1_255(
      {stage09[45]},
      {stage09[63]}
   );
   gpc207_4 gpc207_4_256(
      {stage09[46], stage09[47], stage09[48], stage09[49], stage09[50], stage09[51], stage09[52]},
      {stage11[32], stage11[33]},
      {stage12[47], stage11[47], stage10[50], stage09[64]}
   );
   gpc1_1 gpc1_1_257(
      {stage10[38]},
      {stage10[51]}
   );
   gpc1_1 gpc1_1_258(
      {stage10[39]},
      {stage10[52]}
   );
   gpc1_1 gpc1_1_259(
      {stage10[40]},
      {stage10[53]}
   );
   gpc1_1 gpc1_1_260(
      {stage10[41]},
      {stage10[54]}
   );
   gpc615_5 gpc615_5_261(
      {stage10[42], stage10[43], stage10[44], stage10[45], stage10[46]},
      {stage11[34]},
      {stage12[32], stage12[33], stage12[34], stage12[35], stage12[36], stage12[37]},
      {stage14[50], stage13[48], stage12[48], stage11[48], stage10[55]}
   );
   gpc615_5 gpc615_5_262(
      {stage11[35], stage11[36], stage11[37], stage11[38], stage11[39]},
      {stage12[38]},
      {stage13[32], stage13[33], stage13[34], stage13[35], stage13[36], stage13[37]},
      {stage15[44], stage14[51], stage13[49], stage12[49], stage11[49]}
   );
   gpc615_5 gpc615_5_263(
      {stage11[40], stage11[41], stage11[42], stage11[43], stage11[44]},
      {stage12[39]},
      {stage13[38], stage13[39], stage13[40], stage13[41], stage13[42], stage13[43]},
      {stage15[45], stage14[52], stage13[50], stage12[50], stage11[50]}
   );
   gpc1_1 gpc1_1_264(
      {stage12[40]},
      {stage12[51]}
   );
   gpc615_5 gpc615_5_265(
      {stage12[41], stage12[42], stage12[43], stage12[44], stage12[45]},
      {stage13[44]},
      {stage14[32], stage14[33], stage14[34], stage14[35], stage14[36], stage14[37]},
      {stage16[50], stage15[46], stage14[53], stage13[51], stage12[52]}
   );
   gpc1_1 gpc1_1_266(
      {stage13[45]},
      {stage13[52]}
   );
   gpc1_1 gpc1_1_267(
      {stage13[46]},
      {stage13[53]}
   );
   gpc1_1 gpc1_1_268(
      {stage13[47]},
      {stage13[54]}
   );
   gpc606_5 gpc606_5_269(
      {stage14[38], stage14[39], stage14[40], stage14[41], stage14[42], stage14[43]},
      {stage16[32], stage16[33], stage16[34], stage16[35], stage16[36], stage16[37]},
      {stage18[44], stage17[45], stage16[51], stage15[47], stage14[54]}
   );
   gpc606_5 gpc606_5_270(
      {stage14[44], stage14[45], stage14[46], stage14[47], stage14[48], stage14[49]},
      {stage16[38], stage16[39], stage16[40], stage16[41], stage16[42], stage16[43]},
      {stage18[45], stage17[46], stage16[52], stage15[48], stage14[55]}
   );
   gpc1_1 gpc1_1_271(
      {stage15[32]},
      {stage15[49]}
   );
   gpc1_1 gpc1_1_272(
      {stage15[33]},
      {stage15[50]}
   );
   gpc615_5 gpc615_5_273(
      {stage15[34], stage15[35], stage15[36], stage15[37], stage15[38]},
      {stage16[44]},
      {stage17[32], stage17[33], stage17[34], stage17[35], stage17[36], stage17[37]},
      {stage19[47], stage18[46], stage17[47], stage16[53], stage15[51]}
   );
   gpc615_5 gpc615_5_274(
      {stage15[39], stage15[40], stage15[41], stage15[42], stage15[43]},
      {stage16[45]},
      {stage17[38], stage17[39], stage17[40], stage17[41], stage17[42], stage17[43]},
      {stage19[48], stage18[47], stage17[48], stage16[54], stage15[52]}
   );
   gpc1_1 gpc1_1_275(
      {stage16[46]},
      {stage16[55]}
   );
   gpc1_1 gpc1_1_276(
      {stage16[47]},
      {stage16[56]}
   );
   gpc1_1 gpc1_1_277(
      {stage16[48]},
      {stage16[57]}
   );
   gpc1_1 gpc1_1_278(
      {stage16[49]},
      {stage16[58]}
   );
   gpc1_1 gpc1_1_279(
      {stage17[44]},
      {stage17[49]}
   );
   gpc606_5 gpc606_5_280(
      {stage18[32], stage18[33], stage18[34], stage18[35], stage18[36], stage18[37]},
      {stage20[32], stage20[33], stage20[34], stage20[35], stage20[36], stage20[37]},
      {stage22[47], stage21[48], stage20[49], stage19[49], stage18[48]}
   );
   gpc606_5 gpc606_5_281(
      {stage18[38], stage18[39], stage18[40], stage18[41], stage18[42], stage18[43]},
      {stage20[38], stage20[39], stage20[40], stage20[41], stage20[42], stage20[43]},
      {stage22[48], stage21[49], stage20[50], stage19[50], stage18[49]}
   );
   gpc1_1 gpc1_1_282(
      {stage19[32]},
      {stage19[51]}
   );
   gpc1_1 gpc1_1_283(
      {stage19[33]},
      {stage19[52]}
   );
   gpc606_5 gpc606_5_284(
      {stage19[34], stage19[35], stage19[36], stage19[37], stage19[38], stage19[39]},
      {stage21[32], stage21[33], stage21[34], stage21[35], stage21[36], stage21[37]},
      {stage23[49], stage22[49], stage21[50], stage20[51], stage19[53]}
   );
   gpc207_4 gpc207_4_285(
      {stage19[40], stage19[41], stage19[42], stage19[43], stage19[44], stage19[45], stage19[46]},
      {stage21[38], stage21[39]},
      {stage22[50], stage21[51], stage20[52], stage19[54]}
   );
   gpc2135_5 gpc2135_5_286(
      {stage20[44], stage20[45], stage20[46], stage20[47], stage20[48]},
      {stage21[40], stage21[41], stage21[42]},
      {stage22[32]},
      {stage23[32], stage23[33]},
      {stage24[50], stage23[50], stage22[51], stage21[52], stage20[53]}
   );
   gpc615_5 gpc615_5_287(
      {stage21[43], stage21[44], stage21[45], stage21[46], stage21[47]},
      {stage22[33]},
      {stage23[34], stage23[35], stage23[36], stage23[37], stage23[38], stage23[39]},
      {stage25[45], stage24[51], stage23[51], stage22[52], stage21[53]}
   );
   gpc1_1 gpc1_1_288(
      {stage22[34]},
      {stage22[53]}
   );
   gpc1415_5 gpc1415_5_289(
      {stage22[35], stage22[36], stage22[37], stage22[38], stage22[39]},
      {stage23[40]},
      {stage24[32], stage24[33], stage24[34], stage24[35]},
      {stage25[32]},
      {stage26[53], stage25[46], stage24[52], stage23[52], stage22[54]}
   );
   gpc207_4 gpc207_4_290(
      {stage22[40], stage22[41], stage22[42], stage22[43], stage22[44], stage22[45], stage22[46]},
      {stage24[36], stage24[37]},
      {stage25[47], stage24[53], stage23[53], stage22[55]}
   );
   gpc2135_5 gpc2135_5_291(
      {stage23[41], stage23[42], stage23[43], stage23[44], stage23[45]},
      {stage24[38], stage24[39], stage24[40]},
      {stage25[33]},
      {stage26[32], stage26[33]},
      {stage27[50], stage26[54], stage25[48], stage24[54], stage23[54]}
   );
   gpc2135_5 gpc2135_5_292(
      {stage23[46], stage23[47], stage23[48], 1'h0, 1'h0},
      {stage24[41], stage24[42], stage24[43]},
      {stage25[34]},
      {stage26[34], stage26[35]},
      {stage27[51], stage26[55], stage25[49], stage24[55], stage23[55]}
   );
   gpc1_1 gpc1_1_293(
      {stage24[44]},
      {stage24[56]}
   );
   gpc615_5 gpc615_5_294(
      {stage24[45], stage24[46], stage24[47], stage24[48], stage24[49]},
      {stage25[35]},
      {stage26[36], stage26[37], stage26[38], stage26[39], stage26[40], stage26[41]},
      {stage28[55], stage27[52], stage26[56], stage25[50], stage24[57]}
   );
   gpc1_1 gpc1_1_295(
      {stage25[36]},
      {stage25[51]}
   );
   gpc1_1 gpc1_1_296(
      {stage25[37]},
      {stage25[52]}
   );
   gpc1_1 gpc1_1_297(
      {stage25[38]},
      {stage25[53]}
   );
   gpc606_5 gpc606_5_298(
      {stage25[39], stage25[40], stage25[41], stage25[42], stage25[43], stage25[44]},
      {stage27[32], stage27[33], stage27[34], stage27[35], stage27[36], stage27[37]},
      {stage29[46], stage28[56], stage27[53], stage26[57], stage25[54]}
   );
   gpc606_5 gpc606_5_299(
      {stage26[42], stage26[43], stage26[44], stage26[45], stage26[46], stage26[47]},
      {stage28[32], stage28[33], stage28[34], stage28[35], stage28[36], stage28[37]},
      {stage30[53], stage29[47], stage28[57], stage27[54], stage26[58]}
   );
   gpc606_5 gpc606_5_300(
      {stage26[48], stage26[49], stage26[50], stage26[51], stage26[52], 1'h0},
      {stage28[38], stage28[39], stage28[40], stage28[41], stage28[42], stage28[43]},
      {stage30[54], stage29[48], stage28[58], stage27[55], stage26[59]}
   );
   gpc1_1 gpc1_1_301(
      {stage27[38]},
      {stage27[56]}
   );
   gpc1_1 gpc1_1_302(
      {stage27[39]},
      {stage27[57]}
   );
   gpc1_1 gpc1_1_303(
      {stage27[40]},
      {stage27[58]}
   );
   gpc1_1 gpc1_1_304(
      {stage27[41]},
      {stage27[59]}
   );
   gpc1_1 gpc1_1_305(
      {stage27[42]},
      {stage27[60]}
   );
   gpc1_1 gpc1_1_306(
      {stage27[43]},
      {stage27[61]}
   );
   gpc1_1 gpc1_1_307(
      {stage27[44]},
      {stage27[62]}
   );
   gpc615_5 gpc615_5_308(
      {stage27[45], stage27[46], stage27[47], stage27[48], stage27[49]},
      {stage28[44]},
      {stage29[32], stage29[33], stage29[34], stage29[35], stage29[36], stage29[37]},
      {stage31[48], stage30[55], stage29[49], stage28[59], stage27[63]}
   );
   gpc615_5 gpc615_5_309(
      {stage28[45], stage28[46], stage28[47], stage28[48], stage28[49]},
      {stage29[38]},
      {stage30[32], stage30[33], stage30[34], stage30[35], stage30[36], stage30[37]},
      {stage32[7], stage31[49], stage30[56], stage29[50], stage28[60]}
   );
   gpc615_5 gpc615_5_310(
      {stage28[50], stage28[51], stage28[52], stage28[53], stage28[54]},
      {stage29[39]},
      {stage30[38], stage30[39], stage30[40], stage30[41], stage30[42], stage30[43]},
      {stage32[8], stage31[50], stage30[57], stage29[51], stage28[61]}
   );
   gpc1_1 gpc1_1_311(
      {stage29[40]},
      {stage29[52]}
   );
   gpc615_5 gpc615_5_312(
      {stage29[41], stage29[42], stage29[43], stage29[44], stage29[45]},
      {stage30[44]},
      {stage31[32], stage31[33], stage31[34], stage31[35], stage31[36], stage31[37]},
      {stage33[4], stage32[9], stage31[51], stage30[58], stage29[53]}
   );
   gpc1_1 gpc1_1_313(
      {stage30[45]},
      {stage30[59]}
   );
   gpc1_1 gpc1_1_314(
      {stage30[46]},
      {stage30[60]}
   );
   gpc606_5 gpc606_5_315(
      {stage30[47], stage30[48], stage30[49], stage30[50], stage30[51], stage30[52]},
      {stage32[0], stage32[1], stage32[2], stage32[3], stage32[4], stage32[5]},
      {stage34[0], stage33[5], stage32[10], stage31[52], stage30[61]}
   );
   gpc1_1 gpc1_1_316(
      {stage31[38]},
      {stage31[53]}
   );
   gpc1_1 gpc1_1_317(
      {stage31[39]},
      {stage31[54]}
   );
   gpc1_1 gpc1_1_318(
      {stage31[40]},
      {stage31[55]}
   );
   gpc1_1 gpc1_1_319(
      {stage31[41]},
      {stage31[56]}
   );
   gpc1_1 gpc1_1_320(
      {stage31[42]},
      {stage31[57]}
   );
   gpc1_1 gpc1_1_321(
      {stage31[43]},
      {stage31[58]}
   );
   gpc1_1 gpc1_1_322(
      {stage31[44]},
      {stage31[59]}
   );
   gpc1_1 gpc1_1_323(
      {stage31[45]},
      {stage31[60]}
   );
   gpc1_1 gpc1_1_324(
      {stage31[46]},
      {stage31[61]}
   );
   gpc1_1 gpc1_1_325(
      {stage31[47]},
      {stage31[62]}
   );
   gpc1_1 gpc1_1_326(
      {stage32[6]},
      {stage32[11]}
   );
   gpc1_1 gpc1_1_327(
      {stage33[0]},
      {stage33[6]}
   );
   gpc1_1 gpc1_1_328(
      {stage33[1]},
      {stage33[7]}
   );
   gpc1_1 gpc1_1_329(
      {stage33[2]},
      {stage33[8]}
   );
   gpc1_1 gpc1_1_330(
      {stage33[3]},
      {stage33[9]}
   );
   gpc1_1 gpc1_1_331(
      {stage00[44]},
      {stage00[48]}
   );
   gpc1343_5 gpc1343_5_332(
      {stage00[45], stage00[46], stage00[47]},
      {stage01[44], stage01[45], stage01[46], stage01[47]},
      {stage02[43], stage02[44], stage02[45]},
      {stage03[49]},
      {stage04[64], stage03[56], stage02[51], stage01[48], stage00[49]}
   );
   gpc1_1 gpc1_1_333(
      {stage02[46]},
      {stage02[52]}
   );
   gpc1_1 gpc1_1_334(
      {stage02[47]},
      {stage02[53]}
   );
   gpc223_4 gpc223_4_335(
      {stage02[48], stage02[49], stage02[50]},
      {stage03[50], stage03[51]},
      {stage04[54], stage04[55]},
      {stage05[57], stage04[65], stage03[57], stage02[54]}
   );
   gpc615_5 gpc615_5_336(
      {stage03[52], stage03[53], stage03[54], stage03[55], 1'h0},
      {stage04[56]},
      {stage05[50], stage05[51], stage05[52], stage05[53], stage05[54], stage05[55]},
      {stage07[56], stage06[48], stage05[58], stage04[66], stage03[58]}
   );
   gpc1_1 gpc1_1_337(
      {stage04[57]},
      {stage04[67]}
   );
   gpc1_1 gpc1_1_338(
      {stage04[58]},
      {stage04[68]}
   );
   gpc615_5 gpc615_5_339(
      {stage04[59], stage04[60], stage04[61], stage04[62], stage04[63]},
      {stage05[56]},
      {stage06[42], stage06[43], stage06[44], stage06[45], stage06[46], stage06[47]},
      {stage08[52], stage07[57], stage06[49], stage05[59], stage04[69]}
   );
   gpc2135_5 gpc2135_5_340(
      {stage07[46], stage07[47], stage07[48], stage07[49], stage07[50]},
      {stage08[46], stage08[47], stage08[48]},
      {stage09[53]},
      {stage10[47], stage10[48]},
      {stage11[51], stage10[56], stage09[65], stage08[53], stage07[58]}
   );
   gpc2135_5 gpc2135_5_341(
      {stage07[51], stage07[52], stage07[53], stage07[54], stage07[55]},
      {stage08[49], stage08[50], stage08[51]},
      {stage09[54]},
      {stage10[49], stage10[50]},
      {stage11[52], stage10[57], stage09[66], stage08[54], stage07[59]}
   );
   gpc615_5 gpc615_5_342(
      {stage09[55], stage09[56], stage09[57], stage09[58], stage09[59]},
      {stage10[51]},
      {stage11[45], stage11[46], stage11[47], stage11[48], stage11[49], stage11[50]},
      {stage13[55], stage12[53], stage11[53], stage10[58], stage09[67]}
   );
   gpc2135_5 gpc2135_5_343(
      {stage09[60], stage09[61], stage09[62], stage09[63], stage09[64]},
      {stage10[52], stage10[53], stage10[54]},
      {1'h0},
      {stage12[46], stage12[47]},
      {stage13[56], stage12[54], stage11[54], stage10[59], stage09[68]}
   );
   gpc1_1 gpc1_1_344(
      {stage10[55]},
      {stage10[60]}
   );
   gpc606_5 gpc606_5_345(
      {stage12[48], stage12[49], stage12[50], stage12[51], stage12[52], 1'h0},
      {stage14[50], stage14[51], stage14[52], stage14[53], stage14[54], stage14[55]},
      {stage16[59], stage15[53], stage14[56], stage13[57], stage12[55]}
   );
   gpc207_4 gpc207_4_346(
      {stage13[48], stage13[49], stage13[50], stage13[51], stage13[52], stage13[53], stage13[54]},
      {stage15[44], stage15[45]},
      {stage16[60], stage15[54], stage14[57], stage13[58]}
   );
   gpc7_3 gpc7_3_347(
      {stage15[46], stage15[47], stage15[48], stage15[49], stage15[50], stage15[51], stage15[52]},
      {stage17[50], stage16[61], stage15[55]}
   );
   gpc1_1 gpc1_1_348(
      {stage16[50]},
      {stage16[62]}
   );
   gpc1_1 gpc1_1_349(
      {stage16[51]},
      {stage16[63]}
   );
   gpc207_4 gpc207_4_350(
      {stage16[52], stage16[53], stage16[54], stage16[55], stage16[56], stage16[57], stage16[58]},
      {stage18[44], stage18[45]},
      {stage19[55], stage18[50], stage17[51], stage16[64]}
   );
   gpc207_4 gpc207_4_351(
      {stage17[45], stage17[46], stage17[47], stage17[48], stage17[49], 1'h0, 1'h0},
      {stage19[47], stage19[48]},
      {stage20[54], stage19[56], stage18[51], stage17[52]}
   );
   gpc1_1 gpc1_1_352(
      {stage18[46]},
      {stage18[52]}
   );
   gpc1_1 gpc1_1_353(
      {stage18[47]},
      {stage18[53]}
   );
   gpc1_1 gpc1_1_354(
      {stage18[48]},
      {stage18[54]}
   );
   gpc1_1 gpc1_1_355(
      {stage18[49]},
      {stage18[55]}
   );
   gpc1_1 gpc1_1_356(
      {stage19[49]},
      {stage19[57]}
   );
   gpc615_5 gpc615_5_357(
      {stage19[50], stage19[51], stage19[52], stage19[53], stage19[54]},
      {stage20[49]},
      {stage21[48], stage21[49], stage21[50], stage21[51], stage21[52], stage21[53]},
      {stage23[56], stage22[56], stage21[54], stage20[55], stage19[58]}
   );
   gpc1406_5 gpc1406_5_358(
      {stage20[50], stage20[51], stage20[52], stage20[53], 1'h0, 1'h0},
      {stage22[47], stage22[48], stage22[49], stage22[50]},
      {stage23[49]},
      {stage24[58], stage23[57], stage22[57], stage21[55], stage20[56]}
   );
   gpc135_4 gpc135_4_359(
      {stage22[51], stage22[52], stage22[53], stage22[54], stage22[55]},
      {stage23[50], stage23[51], stage23[52]},
      {stage24[50]},
      {stage25[55], stage24[59], stage23[58], stage22[58]}
   );
   gpc1_1 gpc1_1_360(
      {stage23[53]},
      {stage23[59]}
   );
   gpc1_1 gpc1_1_361(
      {stage23[54]},
      {stage23[60]}
   );
   gpc1_1 gpc1_1_362(
      {stage23[55]},
      {stage23[61]}
   );
   gpc207_4 gpc207_4_363(
      {stage24[51], stage24[52], stage24[53], stage24[54], stage24[55], stage24[56], stage24[57]},
      {stage26[53], stage26[54]},
      {stage27[64], stage26[60], stage25[56], stage24[60]}
   );
   gpc615_5 gpc615_5_364(
      {stage25[45], stage25[46], stage25[47], stage25[48], stage25[49]},
      {stage26[55]},
      {stage27[50], stage27[51], stage27[52], stage27[53], stage27[54], stage27[55]},
      {stage29[54], stage28[62], stage27[65], stage26[61], stage25[57]}
   );
   gpc615_5 gpc615_5_365(
      {stage25[50], stage25[51], stage25[52], stage25[53], stage25[54]},
      {stage26[56]},
      {stage27[56], stage27[57], stage27[58], stage27[59], stage27[60], stage27[61]},
      {stage29[55], stage28[63], stage27[66], stage26[62], stage25[58]}
   );
   gpc1_1 gpc1_1_366(
      {stage26[57]},
      {stage26[63]}
   );
   gpc1_1 gpc1_1_367(
      {stage26[58]},
      {stage26[64]}
   );
   gpc1_1 gpc1_1_368(
      {stage26[59]},
      {stage26[65]}
   );
   gpc1_1 gpc1_1_369(
      {stage27[62]},
      {stage27[67]}
   );
   gpc1_1 gpc1_1_370(
      {stage27[63]},
      {stage27[68]}
   );
   gpc207_4 gpc207_4_371(
      {stage28[55], stage28[56], stage28[57], stage28[58], stage28[59], stage28[60], stage28[61]},
      {stage30[53], stage30[54]},
      {stage31[63], stage30[62], stage29[56], stage28[64]}
   );
   gpc1_1 gpc1_1_372(
      {stage29[46]},
      {stage29[57]}
   );
   gpc1_1 gpc1_1_373(
      {stage29[47]},
      {stage29[58]}
   );
   gpc606_5 gpc606_5_374(
      {stage29[48], stage29[49], stage29[50], stage29[51], stage29[52], stage29[53]},
      {stage31[48], stage31[49], stage31[50], stage31[51], stage31[52], stage31[53]},
      {stage33[10], stage32[12], stage31[64], stage30[63], stage29[59]}
   );
   gpc7_3 gpc7_3_375(
      {stage30[55], stage30[56], stage30[57], stage30[58], stage30[59], stage30[60], stage30[61]},
      {stage32[13], stage31[65], stage30[64]}
   );
   gpc1_1 gpc1_1_376(
      {stage31[54]},
      {stage31[66]}
   );
   gpc1415_5 gpc1415_5_377(
      {stage31[55], stage31[56], stage31[57], stage31[58], stage31[59]},
      {stage32[7]},
      {stage33[4], stage33[5], stage33[6], stage33[7]},
      {stage34[0]},
      {stage35[0], stage34[1], stage33[11], stage32[14], stage31[67]}
   );
   gpc1343_5 gpc1343_5_378(
      {stage31[60], stage31[61], stage31[62]},
      {stage32[8], stage32[9], stage32[10], stage32[11]},
      {stage33[8], stage33[9], 1'h0},
      {1'h0},
      {stage35[1], stage34[2], stage33[12], stage32[15], stage31[68]}
   );
   gpc1_1 gpc1_1_379(
      {stage00[48]},
      {stage00[50]}
   );
   gpc1_1 gpc1_1_380(
      {stage00[49]},
      {stage00[51]}
   );
   gpc1_1 gpc1_1_381(
      {stage01[48]},
      {stage01[49]}
   );
   gpc1_1 gpc1_1_382(
      {stage02[51]},
      {stage02[55]}
   );
   gpc623_5 gpc623_5_383(
      {stage02[52], stage02[53], stage02[54]},
      {stage03[56], stage03[57]},
      {stage04[64], stage04[65], stage04[66], stage04[67], stage04[68], stage04[69]},
      {stage06[50], stage05[60], stage04[70], stage03[59], stage02[56]}
   );
   gpc1_1 gpc1_1_384(
      {stage03[58]},
      {stage03[60]}
   );
   gpc23_3 gpc23_3_385(
      {stage05[57], stage05[58], stage05[59]},
      {stage06[48], stage06[49]},
      {stage07[60], stage06[51], stage05[61]}
   );
   gpc215_4 gpc215_4_386(
      {stage07[56], stage07[57], stage07[58], stage07[59], 1'h0},
      {stage08[52]},
      {stage09[65], stage09[66]},
      {stage10[61], stage09[69], stage08[55], stage07[61]}
   );
   gpc623_5 gpc623_5_387(
      {stage08[53], stage08[54], 1'h0},
      {stage09[67], stage09[68]},
      {stage10[56], stage10[57], stage10[58], stage10[59], stage10[60], 1'h0},
      {stage12[56], stage11[55], stage10[62], stage09[70], stage08[56]}
   );
   gpc2135_5 gpc2135_5_388(
      {stage11[51], stage11[52], stage11[53], stage11[54], 1'h0},
      {stage12[53], stage12[54], stage12[55]},
      {stage13[55]},
      {stage14[56], stage14[57]},
      {stage15[56], stage14[58], stage13[59], stage12[57], stage11[56]}
   );
   gpc3_2 gpc3_2_389(
      {stage13[56], stage13[57], stage13[58]},
      {stage14[59], stage13[60]}
   );
   gpc215_4 gpc215_4_390(
      {stage15[53], stage15[54], stage15[55], 1'h0, 1'h0},
      {stage16[59]},
      {stage17[50], stage17[51]},
      {stage18[56], stage17[53], stage16[65], stage15[57]}
   );
   gpc615_5 gpc615_5_391(
      {stage16[60], stage16[61], stage16[62], stage16[63], stage16[64]},
      {stage17[52]},
      {stage18[50], stage18[51], stage18[52], stage18[53], stage18[54], stage18[55]},
      {stage20[57], stage19[59], stage18[57], stage17[54], stage16[66]}
   );
   gpc2135_5 gpc2135_5_392(
      {stage19[55], stage19[56], stage19[57], stage19[58], 1'h0},
      {stage20[54], stage20[55], stage20[56]},
      {stage21[54]},
      {stage22[56], stage22[57]},
      {stage23[62], stage22[59], stage21[56], stage20[58], stage19[60]}
   );
   gpc1_1 gpc1_1_393(
      {stage21[55]},
      {stage21[57]}
   );
   gpc1_1 gpc1_1_394(
      {stage22[58]},
      {stage22[60]}
   );
   gpc207_4 gpc207_4_395(
      {stage23[56], stage23[57], stage23[58], stage23[59], stage23[60], stage23[61], 1'h0},
      {stage25[55], stage25[56]},
      {stage26[66], stage25[59], stage24[61], stage23[63]}
   );
   gpc623_5 gpc623_5_396(
      {stage24[58], stage24[59], stage24[60]},
      {stage25[57], stage25[58]},
      {stage26[60], stage26[61], stage26[62], stage26[63], stage26[64], stage26[65]},
      {stage28[65], stage27[69], stage26[67], stage25[60], stage24[62]}
   );
   gpc2135_5 gpc2135_5_397(
      {stage27[64], stage27[65], stage27[66], stage27[67], stage27[68]},
      {stage28[62], stage28[63], stage28[64]},
      {stage29[54]},
      {stage30[62], stage30[63]},
      {stage31[69], stage30[65], stage29[60], stage28[66], stage27[70]}
   );
   gpc615_5 gpc615_5_398(
      {stage29[55], stage29[56], stage29[57], stage29[58], stage29[59]},
      {stage30[64]},
      {stage31[63], stage31[64], stage31[65], stage31[66], stage31[67], stage31[68]},
      {stage33[13], stage32[16], stage31[70], stage30[66], stage29[61]}
   );
   gpc2135_5 gpc2135_5_399(
      {stage32[12], stage32[13], stage32[14], stage32[15], 1'h0},
      {stage33[10], stage33[11], stage33[12]},
      {stage34[1]},
      {stage35[0], stage35[1]},
      {stage36[0], stage35[2], stage34[3], stage33[14], stage32[17]}
   );
   gpc1_1 gpc1_1_400(
      {stage34[2]},
      {stage34[4]}
   );
endmodule

module behavioral_tester();
   reg [31:0] src00;
   reg [31:0] src01;
   reg [31:0] src02;
   reg [31:0] src03;
   reg [31:0] src04;
   reg [31:0] src05;
   reg [31:0] src06;
   reg [31:0] src07;
   reg [31:0] src08;
   reg [31:0] src09;
   reg [31:0] src10;
   reg [31:0] src11;
   reg [31:0] src12;
   reg [31:0] src13;
   reg [31:0] src14;
   reg [31:0] src15;
   reg [31:0] src16;
   reg [31:0] src17;
   reg [31:0] src18;
   reg [31:0] src19;
   reg [31:0] src20;
   reg [31:0] src21;
   reg [31:0] src22;
   reg [31:0] src23;
   reg [31:0] src24;
   reg [31:0] src25;
   reg [31:0] src26;
   reg [31:0] src27;
   reg [31:0] src28;
   reg [31:0] src29;
   reg [31:0] src30;
   reg [31:0] src31;
   wire [1:0] dst00;
   wire [0:0] dst01;
   wire [1:0] dst02;
   wire [1:0] dst03;
   wire [0:0] dst04;
   wire [1:0] dst05;
   wire [1:0] dst06;
   wire [1:0] dst07;
   wire [1:0] dst08;
   wire [1:0] dst09;
   wire [1:0] dst10;
   wire [1:0] dst11;
   wire [1:0] dst12;
   wire [1:0] dst13;
   wire [1:0] dst14;
   wire [1:0] dst15;
   wire [1:0] dst16;
   wire [1:0] dst17;
   wire [1:0] dst18;
   wire [1:0] dst19;
   wire [1:0] dst20;
   wire [1:0] dst21;
   wire [1:0] dst22;
   wire [1:0] dst23;
   wire [1:0] dst24;
   wire [1:0] dst25;
   wire [1:0] dst26;
   wire [1:0] dst27;
   wire [1:0] dst28;
   wire [1:0] dst29;
   wire [1:0] dst30;
   wire [1:0] dst31;
   wire [1:0] dst32;
   wire [1:0] dst33;
   wire [1:0] dst34;
   wire [0:0] dst35;
   wire [0:0] dst36;
   wire [37:0] srcsum;
   wire [37:0] dstsum;
   wire test;
   assign srcsum =
      (src00[0] << 0) +
      (src00[1] << 0) +
      (src00[2] << 0) +
      (src00[3] << 0) +
      (src00[4] << 0) +
      (src00[5] << 0) +
      (src00[6] << 0) +
      (src00[7] << 0) +
      (src00[8] << 0) +
      (src00[9] << 0) +
      (src00[10] << 0) +
      (src00[11] << 0) +
      (src00[12] << 0) +
      (src00[13] << 0) +
      (src00[14] << 0) +
      (src00[15] << 0) +
      (src00[16] << 0) +
      (src00[17] << 0) +
      (src00[18] << 0) +
      (src00[19] << 0) +
      (src00[20] << 0) +
      (src00[21] << 0) +
      (src00[22] << 0) +
      (src00[23] << 0) +
      (src00[24] << 0) +
      (src00[25] << 0) +
      (src00[26] << 0) +
      (src00[27] << 0) +
      (src00[28] << 0) +
      (src00[29] << 0) +
      (src00[30] << 0) +
      (src00[31] << 0) +
      (src01[0] << 1) +
      (src01[1] << 1) +
      (src01[2] << 1) +
      (src01[3] << 1) +
      (src01[4] << 1) +
      (src01[5] << 1) +
      (src01[6] << 1) +
      (src01[7] << 1) +
      (src01[8] << 1) +
      (src01[9] << 1) +
      (src01[10] << 1) +
      (src01[11] << 1) +
      (src01[12] << 1) +
      (src01[13] << 1) +
      (src01[14] << 1) +
      (src01[15] << 1) +
      (src01[16] << 1) +
      (src01[17] << 1) +
      (src01[18] << 1) +
      (src01[19] << 1) +
      (src01[20] << 1) +
      (src01[21] << 1) +
      (src01[22] << 1) +
      (src01[23] << 1) +
      (src01[24] << 1) +
      (src01[25] << 1) +
      (src01[26] << 1) +
      (src01[27] << 1) +
      (src01[28] << 1) +
      (src01[29] << 1) +
      (src01[30] << 1) +
      (src01[31] << 1) +
      (src02[0] << 2) +
      (src02[1] << 2) +
      (src02[2] << 2) +
      (src02[3] << 2) +
      (src02[4] << 2) +
      (src02[5] << 2) +
      (src02[6] << 2) +
      (src02[7] << 2) +
      (src02[8] << 2) +
      (src02[9] << 2) +
      (src02[10] << 2) +
      (src02[11] << 2) +
      (src02[12] << 2) +
      (src02[13] << 2) +
      (src02[14] << 2) +
      (src02[15] << 2) +
      (src02[16] << 2) +
      (src02[17] << 2) +
      (src02[18] << 2) +
      (src02[19] << 2) +
      (src02[20] << 2) +
      (src02[21] << 2) +
      (src02[22] << 2) +
      (src02[23] << 2) +
      (src02[24] << 2) +
      (src02[25] << 2) +
      (src02[26] << 2) +
      (src02[27] << 2) +
      (src02[28] << 2) +
      (src02[29] << 2) +
      (src02[30] << 2) +
      (src02[31] << 2) +
      (src03[0] << 3) +
      (src03[1] << 3) +
      (src03[2] << 3) +
      (src03[3] << 3) +
      (src03[4] << 3) +
      (src03[5] << 3) +
      (src03[6] << 3) +
      (src03[7] << 3) +
      (src03[8] << 3) +
      (src03[9] << 3) +
      (src03[10] << 3) +
      (src03[11] << 3) +
      (src03[12] << 3) +
      (src03[13] << 3) +
      (src03[14] << 3) +
      (src03[15] << 3) +
      (src03[16] << 3) +
      (src03[17] << 3) +
      (src03[18] << 3) +
      (src03[19] << 3) +
      (src03[20] << 3) +
      (src03[21] << 3) +
      (src03[22] << 3) +
      (src03[23] << 3) +
      (src03[24] << 3) +
      (src03[25] << 3) +
      (src03[26] << 3) +
      (src03[27] << 3) +
      (src03[28] << 3) +
      (src03[29] << 3) +
      (src03[30] << 3) +
      (src03[31] << 3) +
      (src04[0] << 4) +
      (src04[1] << 4) +
      (src04[2] << 4) +
      (src04[3] << 4) +
      (src04[4] << 4) +
      (src04[5] << 4) +
      (src04[6] << 4) +
      (src04[7] << 4) +
      (src04[8] << 4) +
      (src04[9] << 4) +
      (src04[10] << 4) +
      (src04[11] << 4) +
      (src04[12] << 4) +
      (src04[13] << 4) +
      (src04[14] << 4) +
      (src04[15] << 4) +
      (src04[16] << 4) +
      (src04[17] << 4) +
      (src04[18] << 4) +
      (src04[19] << 4) +
      (src04[20] << 4) +
      (src04[21] << 4) +
      (src04[22] << 4) +
      (src04[23] << 4) +
      (src04[24] << 4) +
      (src04[25] << 4) +
      (src04[26] << 4) +
      (src04[27] << 4) +
      (src04[28] << 4) +
      (src04[29] << 4) +
      (src04[30] << 4) +
      (src04[31] << 4) +
      (src05[0] << 5) +
      (src05[1] << 5) +
      (src05[2] << 5) +
      (src05[3] << 5) +
      (src05[4] << 5) +
      (src05[5] << 5) +
      (src05[6] << 5) +
      (src05[7] << 5) +
      (src05[8] << 5) +
      (src05[9] << 5) +
      (src05[10] << 5) +
      (src05[11] << 5) +
      (src05[12] << 5) +
      (src05[13] << 5) +
      (src05[14] << 5) +
      (src05[15] << 5) +
      (src05[16] << 5) +
      (src05[17] << 5) +
      (src05[18] << 5) +
      (src05[19] << 5) +
      (src05[20] << 5) +
      (src05[21] << 5) +
      (src05[22] << 5) +
      (src05[23] << 5) +
      (src05[24] << 5) +
      (src05[25] << 5) +
      (src05[26] << 5) +
      (src05[27] << 5) +
      (src05[28] << 5) +
      (src05[29] << 5) +
      (src05[30] << 5) +
      (src05[31] << 5) +
      (src06[0] << 6) +
      (src06[1] << 6) +
      (src06[2] << 6) +
      (src06[3] << 6) +
      (src06[4] << 6) +
      (src06[5] << 6) +
      (src06[6] << 6) +
      (src06[7] << 6) +
      (src06[8] << 6) +
      (src06[9] << 6) +
      (src06[10] << 6) +
      (src06[11] << 6) +
      (src06[12] << 6) +
      (src06[13] << 6) +
      (src06[14] << 6) +
      (src06[15] << 6) +
      (src06[16] << 6) +
      (src06[17] << 6) +
      (src06[18] << 6) +
      (src06[19] << 6) +
      (src06[20] << 6) +
      (src06[21] << 6) +
      (src06[22] << 6) +
      (src06[23] << 6) +
      (src06[24] << 6) +
      (src06[25] << 6) +
      (src06[26] << 6) +
      (src06[27] << 6) +
      (src06[28] << 6) +
      (src06[29] << 6) +
      (src06[30] << 6) +
      (src06[31] << 6) +
      (src07[0] << 7) +
      (src07[1] << 7) +
      (src07[2] << 7) +
      (src07[3] << 7) +
      (src07[4] << 7) +
      (src07[5] << 7) +
      (src07[6] << 7) +
      (src07[7] << 7) +
      (src07[8] << 7) +
      (src07[9] << 7) +
      (src07[10] << 7) +
      (src07[11] << 7) +
      (src07[12] << 7) +
      (src07[13] << 7) +
      (src07[14] << 7) +
      (src07[15] << 7) +
      (src07[16] << 7) +
      (src07[17] << 7) +
      (src07[18] << 7) +
      (src07[19] << 7) +
      (src07[20] << 7) +
      (src07[21] << 7) +
      (src07[22] << 7) +
      (src07[23] << 7) +
      (src07[24] << 7) +
      (src07[25] << 7) +
      (src07[26] << 7) +
      (src07[27] << 7) +
      (src07[28] << 7) +
      (src07[29] << 7) +
      (src07[30] << 7) +
      (src07[31] << 7) +
      (src08[0] << 8) +
      (src08[1] << 8) +
      (src08[2] << 8) +
      (src08[3] << 8) +
      (src08[4] << 8) +
      (src08[5] << 8) +
      (src08[6] << 8) +
      (src08[7] << 8) +
      (src08[8] << 8) +
      (src08[9] << 8) +
      (src08[10] << 8) +
      (src08[11] << 8) +
      (src08[12] << 8) +
      (src08[13] << 8) +
      (src08[14] << 8) +
      (src08[15] << 8) +
      (src08[16] << 8) +
      (src08[17] << 8) +
      (src08[18] << 8) +
      (src08[19] << 8) +
      (src08[20] << 8) +
      (src08[21] << 8) +
      (src08[22] << 8) +
      (src08[23] << 8) +
      (src08[24] << 8) +
      (src08[25] << 8) +
      (src08[26] << 8) +
      (src08[27] << 8) +
      (src08[28] << 8) +
      (src08[29] << 8) +
      (src08[30] << 8) +
      (src08[31] << 8) +
      (src09[0] << 9) +
      (src09[1] << 9) +
      (src09[2] << 9) +
      (src09[3] << 9) +
      (src09[4] << 9) +
      (src09[5] << 9) +
      (src09[6] << 9) +
      (src09[7] << 9) +
      (src09[8] << 9) +
      (src09[9] << 9) +
      (src09[10] << 9) +
      (src09[11] << 9) +
      (src09[12] << 9) +
      (src09[13] << 9) +
      (src09[14] << 9) +
      (src09[15] << 9) +
      (src09[16] << 9) +
      (src09[17] << 9) +
      (src09[18] << 9) +
      (src09[19] << 9) +
      (src09[20] << 9) +
      (src09[21] << 9) +
      (src09[22] << 9) +
      (src09[23] << 9) +
      (src09[24] << 9) +
      (src09[25] << 9) +
      (src09[26] << 9) +
      (src09[27] << 9) +
      (src09[28] << 9) +
      (src09[29] << 9) +
      (src09[30] << 9) +
      (src09[31] << 9) +
      (src10[0] << 10) +
      (src10[1] << 10) +
      (src10[2] << 10) +
      (src10[3] << 10) +
      (src10[4] << 10) +
      (src10[5] << 10) +
      (src10[6] << 10) +
      (src10[7] << 10) +
      (src10[8] << 10) +
      (src10[9] << 10) +
      (src10[10] << 10) +
      (src10[11] << 10) +
      (src10[12] << 10) +
      (src10[13] << 10) +
      (src10[14] << 10) +
      (src10[15] << 10) +
      (src10[16] << 10) +
      (src10[17] << 10) +
      (src10[18] << 10) +
      (src10[19] << 10) +
      (src10[20] << 10) +
      (src10[21] << 10) +
      (src10[22] << 10) +
      (src10[23] << 10) +
      (src10[24] << 10) +
      (src10[25] << 10) +
      (src10[26] << 10) +
      (src10[27] << 10) +
      (src10[28] << 10) +
      (src10[29] << 10) +
      (src10[30] << 10) +
      (src10[31] << 10) +
      (src11[0] << 11) +
      (src11[1] << 11) +
      (src11[2] << 11) +
      (src11[3] << 11) +
      (src11[4] << 11) +
      (src11[5] << 11) +
      (src11[6] << 11) +
      (src11[7] << 11) +
      (src11[8] << 11) +
      (src11[9] << 11) +
      (src11[10] << 11) +
      (src11[11] << 11) +
      (src11[12] << 11) +
      (src11[13] << 11) +
      (src11[14] << 11) +
      (src11[15] << 11) +
      (src11[16] << 11) +
      (src11[17] << 11) +
      (src11[18] << 11) +
      (src11[19] << 11) +
      (src11[20] << 11) +
      (src11[21] << 11) +
      (src11[22] << 11) +
      (src11[23] << 11) +
      (src11[24] << 11) +
      (src11[25] << 11) +
      (src11[26] << 11) +
      (src11[27] << 11) +
      (src11[28] << 11) +
      (src11[29] << 11) +
      (src11[30] << 11) +
      (src11[31] << 11) +
      (src12[0] << 12) +
      (src12[1] << 12) +
      (src12[2] << 12) +
      (src12[3] << 12) +
      (src12[4] << 12) +
      (src12[5] << 12) +
      (src12[6] << 12) +
      (src12[7] << 12) +
      (src12[8] << 12) +
      (src12[9] << 12) +
      (src12[10] << 12) +
      (src12[11] << 12) +
      (src12[12] << 12) +
      (src12[13] << 12) +
      (src12[14] << 12) +
      (src12[15] << 12) +
      (src12[16] << 12) +
      (src12[17] << 12) +
      (src12[18] << 12) +
      (src12[19] << 12) +
      (src12[20] << 12) +
      (src12[21] << 12) +
      (src12[22] << 12) +
      (src12[23] << 12) +
      (src12[24] << 12) +
      (src12[25] << 12) +
      (src12[26] << 12) +
      (src12[27] << 12) +
      (src12[28] << 12) +
      (src12[29] << 12) +
      (src12[30] << 12) +
      (src12[31] << 12) +
      (src13[0] << 13) +
      (src13[1] << 13) +
      (src13[2] << 13) +
      (src13[3] << 13) +
      (src13[4] << 13) +
      (src13[5] << 13) +
      (src13[6] << 13) +
      (src13[7] << 13) +
      (src13[8] << 13) +
      (src13[9] << 13) +
      (src13[10] << 13) +
      (src13[11] << 13) +
      (src13[12] << 13) +
      (src13[13] << 13) +
      (src13[14] << 13) +
      (src13[15] << 13) +
      (src13[16] << 13) +
      (src13[17] << 13) +
      (src13[18] << 13) +
      (src13[19] << 13) +
      (src13[20] << 13) +
      (src13[21] << 13) +
      (src13[22] << 13) +
      (src13[23] << 13) +
      (src13[24] << 13) +
      (src13[25] << 13) +
      (src13[26] << 13) +
      (src13[27] << 13) +
      (src13[28] << 13) +
      (src13[29] << 13) +
      (src13[30] << 13) +
      (src13[31] << 13) +
      (src14[0] << 14) +
      (src14[1] << 14) +
      (src14[2] << 14) +
      (src14[3] << 14) +
      (src14[4] << 14) +
      (src14[5] << 14) +
      (src14[6] << 14) +
      (src14[7] << 14) +
      (src14[8] << 14) +
      (src14[9] << 14) +
      (src14[10] << 14) +
      (src14[11] << 14) +
      (src14[12] << 14) +
      (src14[13] << 14) +
      (src14[14] << 14) +
      (src14[15] << 14) +
      (src14[16] << 14) +
      (src14[17] << 14) +
      (src14[18] << 14) +
      (src14[19] << 14) +
      (src14[20] << 14) +
      (src14[21] << 14) +
      (src14[22] << 14) +
      (src14[23] << 14) +
      (src14[24] << 14) +
      (src14[25] << 14) +
      (src14[26] << 14) +
      (src14[27] << 14) +
      (src14[28] << 14) +
      (src14[29] << 14) +
      (src14[30] << 14) +
      (src14[31] << 14) +
      (src15[0] << 15) +
      (src15[1] << 15) +
      (src15[2] << 15) +
      (src15[3] << 15) +
      (src15[4] << 15) +
      (src15[5] << 15) +
      (src15[6] << 15) +
      (src15[7] << 15) +
      (src15[8] << 15) +
      (src15[9] << 15) +
      (src15[10] << 15) +
      (src15[11] << 15) +
      (src15[12] << 15) +
      (src15[13] << 15) +
      (src15[14] << 15) +
      (src15[15] << 15) +
      (src15[16] << 15) +
      (src15[17] << 15) +
      (src15[18] << 15) +
      (src15[19] << 15) +
      (src15[20] << 15) +
      (src15[21] << 15) +
      (src15[22] << 15) +
      (src15[23] << 15) +
      (src15[24] << 15) +
      (src15[25] << 15) +
      (src15[26] << 15) +
      (src15[27] << 15) +
      (src15[28] << 15) +
      (src15[29] << 15) +
      (src15[30] << 15) +
      (src15[31] << 15) +
      (src16[0] << 16) +
      (src16[1] << 16) +
      (src16[2] << 16) +
      (src16[3] << 16) +
      (src16[4] << 16) +
      (src16[5] << 16) +
      (src16[6] << 16) +
      (src16[7] << 16) +
      (src16[8] << 16) +
      (src16[9] << 16) +
      (src16[10] << 16) +
      (src16[11] << 16) +
      (src16[12] << 16) +
      (src16[13] << 16) +
      (src16[14] << 16) +
      (src16[15] << 16) +
      (src16[16] << 16) +
      (src16[17] << 16) +
      (src16[18] << 16) +
      (src16[19] << 16) +
      (src16[20] << 16) +
      (src16[21] << 16) +
      (src16[22] << 16) +
      (src16[23] << 16) +
      (src16[24] << 16) +
      (src16[25] << 16) +
      (src16[26] << 16) +
      (src16[27] << 16) +
      (src16[28] << 16) +
      (src16[29] << 16) +
      (src16[30] << 16) +
      (src16[31] << 16) +
      (src17[0] << 17) +
      (src17[1] << 17) +
      (src17[2] << 17) +
      (src17[3] << 17) +
      (src17[4] << 17) +
      (src17[5] << 17) +
      (src17[6] << 17) +
      (src17[7] << 17) +
      (src17[8] << 17) +
      (src17[9] << 17) +
      (src17[10] << 17) +
      (src17[11] << 17) +
      (src17[12] << 17) +
      (src17[13] << 17) +
      (src17[14] << 17) +
      (src17[15] << 17) +
      (src17[16] << 17) +
      (src17[17] << 17) +
      (src17[18] << 17) +
      (src17[19] << 17) +
      (src17[20] << 17) +
      (src17[21] << 17) +
      (src17[22] << 17) +
      (src17[23] << 17) +
      (src17[24] << 17) +
      (src17[25] << 17) +
      (src17[26] << 17) +
      (src17[27] << 17) +
      (src17[28] << 17) +
      (src17[29] << 17) +
      (src17[30] << 17) +
      (src17[31] << 17) +
      (src18[0] << 18) +
      (src18[1] << 18) +
      (src18[2] << 18) +
      (src18[3] << 18) +
      (src18[4] << 18) +
      (src18[5] << 18) +
      (src18[6] << 18) +
      (src18[7] << 18) +
      (src18[8] << 18) +
      (src18[9] << 18) +
      (src18[10] << 18) +
      (src18[11] << 18) +
      (src18[12] << 18) +
      (src18[13] << 18) +
      (src18[14] << 18) +
      (src18[15] << 18) +
      (src18[16] << 18) +
      (src18[17] << 18) +
      (src18[18] << 18) +
      (src18[19] << 18) +
      (src18[20] << 18) +
      (src18[21] << 18) +
      (src18[22] << 18) +
      (src18[23] << 18) +
      (src18[24] << 18) +
      (src18[25] << 18) +
      (src18[26] << 18) +
      (src18[27] << 18) +
      (src18[28] << 18) +
      (src18[29] << 18) +
      (src18[30] << 18) +
      (src18[31] << 18) +
      (src19[0] << 19) +
      (src19[1] << 19) +
      (src19[2] << 19) +
      (src19[3] << 19) +
      (src19[4] << 19) +
      (src19[5] << 19) +
      (src19[6] << 19) +
      (src19[7] << 19) +
      (src19[8] << 19) +
      (src19[9] << 19) +
      (src19[10] << 19) +
      (src19[11] << 19) +
      (src19[12] << 19) +
      (src19[13] << 19) +
      (src19[14] << 19) +
      (src19[15] << 19) +
      (src19[16] << 19) +
      (src19[17] << 19) +
      (src19[18] << 19) +
      (src19[19] << 19) +
      (src19[20] << 19) +
      (src19[21] << 19) +
      (src19[22] << 19) +
      (src19[23] << 19) +
      (src19[24] << 19) +
      (src19[25] << 19) +
      (src19[26] << 19) +
      (src19[27] << 19) +
      (src19[28] << 19) +
      (src19[29] << 19) +
      (src19[30] << 19) +
      (src19[31] << 19) +
      (src20[0] << 20) +
      (src20[1] << 20) +
      (src20[2] << 20) +
      (src20[3] << 20) +
      (src20[4] << 20) +
      (src20[5] << 20) +
      (src20[6] << 20) +
      (src20[7] << 20) +
      (src20[8] << 20) +
      (src20[9] << 20) +
      (src20[10] << 20) +
      (src20[11] << 20) +
      (src20[12] << 20) +
      (src20[13] << 20) +
      (src20[14] << 20) +
      (src20[15] << 20) +
      (src20[16] << 20) +
      (src20[17] << 20) +
      (src20[18] << 20) +
      (src20[19] << 20) +
      (src20[20] << 20) +
      (src20[21] << 20) +
      (src20[22] << 20) +
      (src20[23] << 20) +
      (src20[24] << 20) +
      (src20[25] << 20) +
      (src20[26] << 20) +
      (src20[27] << 20) +
      (src20[28] << 20) +
      (src20[29] << 20) +
      (src20[30] << 20) +
      (src20[31] << 20) +
      (src21[0] << 21) +
      (src21[1] << 21) +
      (src21[2] << 21) +
      (src21[3] << 21) +
      (src21[4] << 21) +
      (src21[5] << 21) +
      (src21[6] << 21) +
      (src21[7] << 21) +
      (src21[8] << 21) +
      (src21[9] << 21) +
      (src21[10] << 21) +
      (src21[11] << 21) +
      (src21[12] << 21) +
      (src21[13] << 21) +
      (src21[14] << 21) +
      (src21[15] << 21) +
      (src21[16] << 21) +
      (src21[17] << 21) +
      (src21[18] << 21) +
      (src21[19] << 21) +
      (src21[20] << 21) +
      (src21[21] << 21) +
      (src21[22] << 21) +
      (src21[23] << 21) +
      (src21[24] << 21) +
      (src21[25] << 21) +
      (src21[26] << 21) +
      (src21[27] << 21) +
      (src21[28] << 21) +
      (src21[29] << 21) +
      (src21[30] << 21) +
      (src21[31] << 21) +
      (src22[0] << 22) +
      (src22[1] << 22) +
      (src22[2] << 22) +
      (src22[3] << 22) +
      (src22[4] << 22) +
      (src22[5] << 22) +
      (src22[6] << 22) +
      (src22[7] << 22) +
      (src22[8] << 22) +
      (src22[9] << 22) +
      (src22[10] << 22) +
      (src22[11] << 22) +
      (src22[12] << 22) +
      (src22[13] << 22) +
      (src22[14] << 22) +
      (src22[15] << 22) +
      (src22[16] << 22) +
      (src22[17] << 22) +
      (src22[18] << 22) +
      (src22[19] << 22) +
      (src22[20] << 22) +
      (src22[21] << 22) +
      (src22[22] << 22) +
      (src22[23] << 22) +
      (src22[24] << 22) +
      (src22[25] << 22) +
      (src22[26] << 22) +
      (src22[27] << 22) +
      (src22[28] << 22) +
      (src22[29] << 22) +
      (src22[30] << 22) +
      (src22[31] << 22) +
      (src23[0] << 23) +
      (src23[1] << 23) +
      (src23[2] << 23) +
      (src23[3] << 23) +
      (src23[4] << 23) +
      (src23[5] << 23) +
      (src23[6] << 23) +
      (src23[7] << 23) +
      (src23[8] << 23) +
      (src23[9] << 23) +
      (src23[10] << 23) +
      (src23[11] << 23) +
      (src23[12] << 23) +
      (src23[13] << 23) +
      (src23[14] << 23) +
      (src23[15] << 23) +
      (src23[16] << 23) +
      (src23[17] << 23) +
      (src23[18] << 23) +
      (src23[19] << 23) +
      (src23[20] << 23) +
      (src23[21] << 23) +
      (src23[22] << 23) +
      (src23[23] << 23) +
      (src23[24] << 23) +
      (src23[25] << 23) +
      (src23[26] << 23) +
      (src23[27] << 23) +
      (src23[28] << 23) +
      (src23[29] << 23) +
      (src23[30] << 23) +
      (src23[31] << 23) +
      (src24[0] << 24) +
      (src24[1] << 24) +
      (src24[2] << 24) +
      (src24[3] << 24) +
      (src24[4] << 24) +
      (src24[5] << 24) +
      (src24[6] << 24) +
      (src24[7] << 24) +
      (src24[8] << 24) +
      (src24[9] << 24) +
      (src24[10] << 24) +
      (src24[11] << 24) +
      (src24[12] << 24) +
      (src24[13] << 24) +
      (src24[14] << 24) +
      (src24[15] << 24) +
      (src24[16] << 24) +
      (src24[17] << 24) +
      (src24[18] << 24) +
      (src24[19] << 24) +
      (src24[20] << 24) +
      (src24[21] << 24) +
      (src24[22] << 24) +
      (src24[23] << 24) +
      (src24[24] << 24) +
      (src24[25] << 24) +
      (src24[26] << 24) +
      (src24[27] << 24) +
      (src24[28] << 24) +
      (src24[29] << 24) +
      (src24[30] << 24) +
      (src24[31] << 24) +
      (src25[0] << 25) +
      (src25[1] << 25) +
      (src25[2] << 25) +
      (src25[3] << 25) +
      (src25[4] << 25) +
      (src25[5] << 25) +
      (src25[6] << 25) +
      (src25[7] << 25) +
      (src25[8] << 25) +
      (src25[9] << 25) +
      (src25[10] << 25) +
      (src25[11] << 25) +
      (src25[12] << 25) +
      (src25[13] << 25) +
      (src25[14] << 25) +
      (src25[15] << 25) +
      (src25[16] << 25) +
      (src25[17] << 25) +
      (src25[18] << 25) +
      (src25[19] << 25) +
      (src25[20] << 25) +
      (src25[21] << 25) +
      (src25[22] << 25) +
      (src25[23] << 25) +
      (src25[24] << 25) +
      (src25[25] << 25) +
      (src25[26] << 25) +
      (src25[27] << 25) +
      (src25[28] << 25) +
      (src25[29] << 25) +
      (src25[30] << 25) +
      (src25[31] << 25) +
      (src26[0] << 26) +
      (src26[1] << 26) +
      (src26[2] << 26) +
      (src26[3] << 26) +
      (src26[4] << 26) +
      (src26[5] << 26) +
      (src26[6] << 26) +
      (src26[7] << 26) +
      (src26[8] << 26) +
      (src26[9] << 26) +
      (src26[10] << 26) +
      (src26[11] << 26) +
      (src26[12] << 26) +
      (src26[13] << 26) +
      (src26[14] << 26) +
      (src26[15] << 26) +
      (src26[16] << 26) +
      (src26[17] << 26) +
      (src26[18] << 26) +
      (src26[19] << 26) +
      (src26[20] << 26) +
      (src26[21] << 26) +
      (src26[22] << 26) +
      (src26[23] << 26) +
      (src26[24] << 26) +
      (src26[25] << 26) +
      (src26[26] << 26) +
      (src26[27] << 26) +
      (src26[28] << 26) +
      (src26[29] << 26) +
      (src26[30] << 26) +
      (src26[31] << 26) +
      (src27[0] << 27) +
      (src27[1] << 27) +
      (src27[2] << 27) +
      (src27[3] << 27) +
      (src27[4] << 27) +
      (src27[5] << 27) +
      (src27[6] << 27) +
      (src27[7] << 27) +
      (src27[8] << 27) +
      (src27[9] << 27) +
      (src27[10] << 27) +
      (src27[11] << 27) +
      (src27[12] << 27) +
      (src27[13] << 27) +
      (src27[14] << 27) +
      (src27[15] << 27) +
      (src27[16] << 27) +
      (src27[17] << 27) +
      (src27[18] << 27) +
      (src27[19] << 27) +
      (src27[20] << 27) +
      (src27[21] << 27) +
      (src27[22] << 27) +
      (src27[23] << 27) +
      (src27[24] << 27) +
      (src27[25] << 27) +
      (src27[26] << 27) +
      (src27[27] << 27) +
      (src27[28] << 27) +
      (src27[29] << 27) +
      (src27[30] << 27) +
      (src27[31] << 27) +
      (src28[0] << 28) +
      (src28[1] << 28) +
      (src28[2] << 28) +
      (src28[3] << 28) +
      (src28[4] << 28) +
      (src28[5] << 28) +
      (src28[6] << 28) +
      (src28[7] << 28) +
      (src28[8] << 28) +
      (src28[9] << 28) +
      (src28[10] << 28) +
      (src28[11] << 28) +
      (src28[12] << 28) +
      (src28[13] << 28) +
      (src28[14] << 28) +
      (src28[15] << 28) +
      (src28[16] << 28) +
      (src28[17] << 28) +
      (src28[18] << 28) +
      (src28[19] << 28) +
      (src28[20] << 28) +
      (src28[21] << 28) +
      (src28[22] << 28) +
      (src28[23] << 28) +
      (src28[24] << 28) +
      (src28[25] << 28) +
      (src28[26] << 28) +
      (src28[27] << 28) +
      (src28[28] << 28) +
      (src28[29] << 28) +
      (src28[30] << 28) +
      (src28[31] << 28) +
      (src29[0] << 29) +
      (src29[1] << 29) +
      (src29[2] << 29) +
      (src29[3] << 29) +
      (src29[4] << 29) +
      (src29[5] << 29) +
      (src29[6] << 29) +
      (src29[7] << 29) +
      (src29[8] << 29) +
      (src29[9] << 29) +
      (src29[10] << 29) +
      (src29[11] << 29) +
      (src29[12] << 29) +
      (src29[13] << 29) +
      (src29[14] << 29) +
      (src29[15] << 29) +
      (src29[16] << 29) +
      (src29[17] << 29) +
      (src29[18] << 29) +
      (src29[19] << 29) +
      (src29[20] << 29) +
      (src29[21] << 29) +
      (src29[22] << 29) +
      (src29[23] << 29) +
      (src29[24] << 29) +
      (src29[25] << 29) +
      (src29[26] << 29) +
      (src29[27] << 29) +
      (src29[28] << 29) +
      (src29[29] << 29) +
      (src29[30] << 29) +
      (src29[31] << 29) +
      (src30[0] << 30) +
      (src30[1] << 30) +
      (src30[2] << 30) +
      (src30[3] << 30) +
      (src30[4] << 30) +
      (src30[5] << 30) +
      (src30[6] << 30) +
      (src30[7] << 30) +
      (src30[8] << 30) +
      (src30[9] << 30) +
      (src30[10] << 30) +
      (src30[11] << 30) +
      (src30[12] << 30) +
      (src30[13] << 30) +
      (src30[14] << 30) +
      (src30[15] << 30) +
      (src30[16] << 30) +
      (src30[17] << 30) +
      (src30[18] << 30) +
      (src30[19] << 30) +
      (src30[20] << 30) +
      (src30[21] << 30) +
      (src30[22] << 30) +
      (src30[23] << 30) +
      (src30[24] << 30) +
      (src30[25] << 30) +
      (src30[26] << 30) +
      (src30[27] << 30) +
      (src30[28] << 30) +
      (src30[29] << 30) +
      (src30[30] << 30) +
      (src30[31] << 30) +
      (src31[0] << 31) +
      (src31[1] << 31) +
      (src31[2] << 31) +
      (src31[3] << 31) +
      (src31[4] << 31) +
      (src31[5] << 31) +
      (src31[6] << 31) +
      (src31[7] << 31) +
      (src31[8] << 31) +
      (src31[9] << 31) +
      (src31[10] << 31) +
      (src31[11] << 31) +
      (src31[12] << 31) +
      (src31[13] << 31) +
      (src31[14] << 31) +
      (src31[15] << 31) +
      (src31[16] << 31) +
      (src31[17] << 31) +
      (src31[18] << 31) +
      (src31[19] << 31) +
      (src31[20] << 31) +
      (src31[21] << 31) +
      (src31[22] << 31) +
      (src31[23] << 31) +
      (src31[24] << 31) +
      (src31[25] << 31) +
      (src31[26] << 31) +
      (src31[27] << 31) +
      (src31[28] << 31) +
      (src31[29] << 31) +
      (src31[30] << 31) +
      (src31[31] << 31);
   assign dstsum =
      (dst00[0] << 0) +
      (dst00[1] << 0) +
      (dst01[0] << 1) +
      (dst02[0] << 2) +
      (dst02[1] << 2) +
      (dst03[0] << 3) +
      (dst03[1] << 3) +
      (dst04[0] << 4) +
      (dst05[0] << 5) +
      (dst05[1] << 5) +
      (dst06[0] << 6) +
      (dst06[1] << 6) +
      (dst07[0] << 7) +
      (dst07[1] << 7) +
      (dst08[0] << 8) +
      (dst08[1] << 8) +
      (dst09[0] << 9) +
      (dst09[1] << 9) +
      (dst10[0] << 10) +
      (dst10[1] << 10) +
      (dst11[0] << 11) +
      (dst11[1] << 11) +
      (dst12[0] << 12) +
      (dst12[1] << 12) +
      (dst13[0] << 13) +
      (dst13[1] << 13) +
      (dst14[0] << 14) +
      (dst14[1] << 14) +
      (dst15[0] << 15) +
      (dst15[1] << 15) +
      (dst16[0] << 16) +
      (dst16[1] << 16) +
      (dst17[0] << 17) +
      (dst17[1] << 17) +
      (dst18[0] << 18) +
      (dst18[1] << 18) +
      (dst19[0] << 19) +
      (dst19[1] << 19) +
      (dst20[0] << 20) +
      (dst20[1] << 20) +
      (dst21[0] << 21) +
      (dst21[1] << 21) +
      (dst22[0] << 22) +
      (dst22[1] << 22) +
      (dst23[0] << 23) +
      (dst23[1] << 23) +
      (dst24[0] << 24) +
      (dst24[1] << 24) +
      (dst25[0] << 25) +
      (dst25[1] << 25) +
      (dst26[0] << 26) +
      (dst26[1] << 26) +
      (dst27[0] << 27) +
      (dst27[1] << 27) +
      (dst28[0] << 28) +
      (dst28[1] << 28) +
      (dst29[0] << 29) +
      (dst29[1] << 29) +
      (dst30[0] << 30) +
      (dst30[1] << 30) +
      (dst31[0] << 31) +
      (dst31[1] << 31) +
      (dst32[0] << 32) +
      (dst32[1] << 32) +
      (dst33[0] << 33) +
      (dst33[1] << 33) +
      (dst34[0] << 34) +
      (dst34[1] << 34) +
      (dst35[0] << 35) +
      (dst36[0] << 36);
   compressor main_cmp(src00, src01, src02, src03, src04, src05, src06, src07, src08, src09, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, dst00, dst01, dst02, dst03, dst04, dst05, dst06, dst07, dst08, dst09, dst10, dst11, dst12, dst13, dst14, dst15, dst16, dst17, dst18, dst19, dst20, dst21, dst22, dst23, dst24, dst25, dst26, dst27, dst28, dst29, dst30, dst31, dst32, dst33, dst34, dst35, dst36);
   assign test = srcsum == dstsum;
   initial begin
      $monitor("src: 0x%x, dst: 0x%x, test: %b", srcsum, dstsum, test);
   end
   initial begin
      src00 <= 32'h0;
      src01 <= 32'h0;
      src02 <= 32'h0;
      src03 <= 32'h0;
      src04 <= 32'h0;
      src05 <= 32'h0;
      src06 <= 32'h0;
      src07 <= 32'h0;
      src08 <= 32'h0;
      src09 <= 32'h0;
      src10 <= 32'h0;
      src11 <= 32'h0;
      src12 <= 32'h0;
      src13 <= 32'h0;
      src14 <= 32'h0;
      src15 <= 32'h0;
      src16 <= 32'h0;
      src17 <= 32'h0;
      src18 <= 32'h0;
      src19 <= 32'h0;
      src20 <= 32'h0;
      src21 <= 32'h0;
      src22 <= 32'h0;
      src23 <= 32'h0;
      src24 <= 32'h0;
      src25 <= 32'h0;
      src26 <= 32'h0;
      src27 <= 32'h0;
      src28 <= 32'h0;
      src29 <= 32'h0;
      src30 <= 32'h0;
      src31 <= 32'h0;
      #1
      src00 <= 32'hffffffff;
      src01 <= 32'hffffffff;
      src02 <= 32'hffffffff;
      src03 <= 32'hffffffff;
      src04 <= 32'hffffffff;
      src05 <= 32'hffffffff;
      src06 <= 32'hffffffff;
      src07 <= 32'hffffffff;
      src08 <= 32'hffffffff;
      src09 <= 32'hffffffff;
      src10 <= 32'hffffffff;
      src11 <= 32'hffffffff;
      src12 <= 32'hffffffff;
      src13 <= 32'hffffffff;
      src14 <= 32'hffffffff;
      src15 <= 32'hffffffff;
      src16 <= 32'hffffffff;
      src17 <= 32'hffffffff;
      src18 <= 32'hffffffff;
      src19 <= 32'hffffffff;
      src20 <= 32'hffffffff;
      src21 <= 32'hffffffff;
      src22 <= 32'hffffffff;
      src23 <= 32'hffffffff;
      src24 <= 32'hffffffff;
      src25 <= 32'hffffffff;
      src26 <= 32'hffffffff;
      src27 <= 32'hffffffff;
      src28 <= 32'hffffffff;
      src29 <= 32'hffffffff;
      src30 <= 32'hffffffff;
      src31 <= 32'hffffffff;
      #1
      src00 <= 32'hd82c07cd;
      src01 <= 32'h6baa9455;
      src02 <= 32'h82e2e662;
      src03 <= 32'h7a024204;
      src04 <= 32'he87a1613;
      src05 <= 32'h81332876;
      src06 <= 32'h48268673;
      src07 <= 32'hc17c6279;
      src08 <= 32'he6f4590b;
      src09 <= 32'h4f65d4d9;
      src10 <= 32'hbad640fb;
      src11 <= 32'haf19922a;
      src12 <= 32'h19c78df4;
      src13 <= 32'h6f25e2a2;
      src14 <= 32'he9bb17bc;
      src15 <= 32'h7a1d5006;
      src16 <= 32'h42af9fc3;
      src17 <= 32'h3983ca8;
      src18 <= 32'hde1b372a;
      src19 <= 32'hded733e8;
      src20 <= 32'h9148624f;
      src21 <= 32'hf7b0b7d2;
      src22 <= 32'h72ae2244;
      src23 <= 32'heece328b;
      src24 <= 32'h1beb3711;
      src25 <= 32'h8d1fd9b7;
      src26 <= 32'hb4e1357d;
      src27 <= 32'h8c25166a;
      src28 <= 32'h8a5006c1;
      src29 <= 32'h966e1277;
      src30 <= 32'h71eacd05;
      src31 <= 32'h6288e1a5;
      #1
      src00 <= 32'h935ddd72;
      src01 <= 32'h4a5308cc;
      src02 <= 32'h2fcd81b5;
      src03 <= 32'ha81ad477;
      src04 <= 32'h79fdef7c;
      src05 <= 32'hc1f254b8;
      src06 <= 32'he07405eb;
      src07 <= 32'hec62b2c8;
      src08 <= 32'hd7ab7928;
      src09 <= 32'hcfc6e625;
      src10 <= 32'hd977e993;
      src11 <= 32'hf323ca74;
      src12 <= 32'h9466e472;
      src13 <= 32'h73581a81;
      src14 <= 32'hcb175a5a;
      src15 <= 32'h15166570;
      src16 <= 32'h9cdf5a86;
      src17 <= 32'ha1515607;
      src18 <= 32'hd8570102;
      src19 <= 32'h3e37952d;
      src20 <= 32'hbb42e0b2;
      src21 <= 32'h38701a14;
      src22 <= 32'hcb69ca38;
      src23 <= 32'h552116dd;
      src24 <= 32'hd0dfae43;
      src25 <= 32'hb29a8b06;
      src26 <= 32'hae3b16ec;
      src27 <= 32'h6d599e8;
      src28 <= 32'ha28f5ab0;
      src29 <= 32'h9371a71f;
      src30 <= 32'h64264cd5;
      src31 <= 32'hfb0323a1;
      #1
      src00 <= 32'h589f877;
      src01 <= 32'h1fb797fa;
      src02 <= 32'hccfdba9b;
      src03 <= 32'h428a1c22;
      src04 <= 32'h38884479;
      src05 <= 32'ha59cec98;
      src06 <= 32'h59acdd98;
      src07 <= 32'h2e295065;
      src08 <= 32'h80ee526e;
      src09 <= 32'hfcfcfa81;
      src10 <= 32'h3308fb2e;
      src11 <= 32'hbb4a06cb;
      src12 <= 32'hac322c12;
      src13 <= 32'had1b8f60;
      src14 <= 32'hd86dbf11;
      src15 <= 32'h402d0baf;
      src16 <= 32'h2cc0f859;
      src17 <= 32'h5b6e4ae7;
      src18 <= 32'h403d1f83;
      src19 <= 32'h32f06ca;
      src20 <= 32'hbdd7d19b;
      src21 <= 32'h47e7f593;
      src22 <= 32'hf40048d7;
      src23 <= 32'h9efee464;
      src24 <= 32'hb732d46f;
      src25 <= 32'ha69cfb85;
      src26 <= 32'h559b5975;
      src27 <= 32'h3d4a5d51;
      src28 <= 32'ha32c9b6f;
      src29 <= 32'h6a1689ad;
      src30 <= 32'hbf9c0ef;
      src31 <= 32'h720299e3;
      #1
      src00 <= 32'h285e25b4;
      src01 <= 32'hc167733f;
      src02 <= 32'he245a460;
      src03 <= 32'h7e9cf84f;
      src04 <= 32'h77863fe5;
      src05 <= 32'hcffa6cdd;
      src06 <= 32'hb9bdee2d;
      src07 <= 32'hfca05536;
      src08 <= 32'hadb328cb;
      src09 <= 32'h50f0fc2b;
      src10 <= 32'h36a98d74;
      src11 <= 32'h19086515;
      src12 <= 32'ha636425c;
      src13 <= 32'hdfa7c6ed;
      src14 <= 32'hfa7ff8bf;
      src15 <= 32'h19a5711b;
      src16 <= 32'h14d30dbc;
      src17 <= 32'hcad6e514;
      src18 <= 32'hdc821527;
      src19 <= 32'h58d87776;
      src20 <= 32'hdf3277fd;
      src21 <= 32'h4c14982;
      src22 <= 32'ha68e88e;
      src23 <= 32'hae55cdff;
      src24 <= 32'h8ef066d4;
      src25 <= 32'hf24dfdd8;
      src26 <= 32'ha7c5cb87;
      src27 <= 32'he7180322;
      src28 <= 32'ha3e04b3b;
      src29 <= 32'h89b5b368;
      src30 <= 32'h35354579;
      src31 <= 32'h964ddb77;
      #1
      src00 <= 32'h247145f;
      src01 <= 32'h26a97465;
      src02 <= 32'h555a4085;
      src03 <= 32'hca24be4d;
      src04 <= 32'hb7ef941c;
      src05 <= 32'h9edb95f2;
      src06 <= 32'ha8c46c7;
      src07 <= 32'h29f2c3c7;
      src08 <= 32'h4a1eb1b7;
      src09 <= 32'h8c69778f;
      src10 <= 32'h4b1cb8bd;
      src11 <= 32'hc5a876f;
      src12 <= 32'h122411e6;
      src13 <= 32'h5419eefc;
      src14 <= 32'h6a2b3200;
      src15 <= 32'he89dc815;
      src16 <= 32'h79585e69;
      src17 <= 32'h57f98d1e;
      src18 <= 32'h7aa56a18;
      src19 <= 32'hb318ad4c;
      src20 <= 32'h6d316b4a;
      src21 <= 32'h4d4985dc;
      src22 <= 32'he4f7625e;
      src23 <= 32'heb70ba65;
      src24 <= 32'ha38d8afc;
      src25 <= 32'h15ace7a1;
      src26 <= 32'hbff773ce;
      src27 <= 32'hfa7ee05;
      src28 <= 32'h202861c;
      src29 <= 32'h84dd6da6;
      src30 <= 32'hade6c5e9;
      src31 <= 32'h6c4c3935;
      #1
      src00 <= 32'h5e4af862;
      src01 <= 32'hc6f00933;
      src02 <= 32'h6e648043;
      src03 <= 32'h5bc7fdeb;
      src04 <= 32'hb3b68b57;
      src05 <= 32'had4ab155;
      src06 <= 32'h1e70e799;
      src07 <= 32'h65e04993;
      src08 <= 32'h25777cf0;
      src09 <= 32'h32ae2a20;
      src10 <= 32'h60c6b3ed;
      src11 <= 32'h26bdd974;
      src12 <= 32'hfba52e59;
      src13 <= 32'hae0fdbc8;
      src14 <= 32'h38018399;
      src15 <= 32'he6256403;
      src16 <= 32'hd17034ce;
      src17 <= 32'hc8bf23fb;
      src18 <= 32'hd7a3283c;
      src19 <= 32'h953c178e;
      src20 <= 32'hce9b2e70;
      src21 <= 32'ha1727f7;
      src22 <= 32'h399f8a8f;
      src23 <= 32'ha66dc4e;
      src24 <= 32'hd80d6a1c;
      src25 <= 32'ha7f5195c;
      src26 <= 32'hf7f60e7f;
      src27 <= 32'h8147a8f4;
      src28 <= 32'h809f2923;
      src29 <= 32'h92e94e89;
      src30 <= 32'hfd938adc;
      src31 <= 32'hbf391fbb;
      #1
      src00 <= 32'h34c3494a;
      src01 <= 32'h993ec8c6;
      src02 <= 32'h961d8dcf;
      src03 <= 32'hcc4da021;
      src04 <= 32'h2e9583ea;
      src05 <= 32'h4124405b;
      src06 <= 32'h10cc8711;
      src07 <= 32'hdc2151e1;
      src08 <= 32'h68777bab;
      src09 <= 32'hcf5e9ea3;
      src10 <= 32'hff030b8;
      src11 <= 32'h209818d1;
      src12 <= 32'hd476fe38;
      src13 <= 32'h932f5b6;
      src14 <= 32'h6af944e0;
      src15 <= 32'hb799ae8e;
      src16 <= 32'hfc98c279;
      src17 <= 32'h69407be7;
      src18 <= 32'h9c9d03f3;
      src19 <= 32'h62fda854;
      src20 <= 32'hc0a5967;
      src21 <= 32'h26c00984;
      src22 <= 32'h9e0df45b;
      src23 <= 32'ha1457899;
      src24 <= 32'h58bf3b9e;
      src25 <= 32'h7d859725;
      src26 <= 32'he19b5837;
      src27 <= 32'h9f3dd894;
      src28 <= 32'he96aa1af;
      src29 <= 32'hcca1a034;
      src30 <= 32'hcf6c9992;
      src31 <= 32'h306aa871;
      #1
      src00 <= 32'hc838a145;
      src01 <= 32'h71cff814;
      src02 <= 32'hc1b199c4;
      src03 <= 32'h7499b28c;
      src04 <= 32'hef2d9a38;
      src05 <= 32'h7c7550f2;
      src06 <= 32'he6ac9d8a;
      src07 <= 32'h374a6cc9;
      src08 <= 32'h1d0ab994;
      src09 <= 32'h90e639e1;
      src10 <= 32'hec41e6f6;
      src11 <= 32'hef8d9ff0;
      src12 <= 32'h6a677623;
      src13 <= 32'h1965e435;
      src14 <= 32'hc618fc1e;
      src15 <= 32'h725c2675;
      src16 <= 32'hafb918c8;
      src17 <= 32'h7b6e08e;
      src18 <= 32'hf655860b;
      src19 <= 32'hb8f8903b;
      src20 <= 32'h141b1a1b;
      src21 <= 32'h12011caa;
      src22 <= 32'h78548d7;
      src23 <= 32'h590e83da;
      src24 <= 32'hf96d4403;
      src25 <= 32'hd1aa6c5e;
      src26 <= 32'he4b82987;
      src27 <= 32'h353e0c86;
      src28 <= 32'h1d6d903;
      src29 <= 32'h9ad7558f;
      src30 <= 32'hdbf2eed1;
      src31 <= 32'h2fdeb035;
      #1
      src00 <= 32'h1cc5a8a0;
      src01 <= 32'hf58c43ce;
      src02 <= 32'h215203c7;
      src03 <= 32'hf76dce6e;
      src04 <= 32'h5cbbc080;
      src05 <= 32'h4ae9ee11;
      src06 <= 32'ha2cb5f38;
      src07 <= 32'hfe3216bd;
      src08 <= 32'h94b28b9d;
      src09 <= 32'h280a07ee;
      src10 <= 32'he5ce0ca6;
      src11 <= 32'hf217faac;
      src12 <= 32'hcdec85da;
      src13 <= 32'h3e2aad3e;
      src14 <= 32'hc13e66af;
      src15 <= 32'h4a82e06a;
      src16 <= 32'h542bd75;
      src17 <= 32'h12bdf75f;
      src18 <= 32'h6b944e09;
      src19 <= 32'h8cffbbb1;
      src20 <= 32'h6c148fc6;
      src21 <= 32'ha31034dd;
      src22 <= 32'h15a5712c;
      src23 <= 32'hecfb95b;
      src24 <= 32'h689bba65;
      src25 <= 32'h52177eb7;
      src26 <= 32'h3438b4e4;
      src27 <= 32'h788c161e;
      src28 <= 32'hf344c911;
      src29 <= 32'hcbe88a3f;
      src30 <= 32'h46e785ad;
      src31 <= 32'hb02de52c;
      #1
      src00 <= 32'h66163e5b;
      src01 <= 32'hc4841a8d;
      src02 <= 32'h6e84f8ea;
      src03 <= 32'h74151acc;
      src04 <= 32'h247f4d97;
      src05 <= 32'ha32652e8;
      src06 <= 32'h3421beaf;
      src07 <= 32'hb2f11ef9;
      src08 <= 32'h9e65736c;
      src09 <= 32'h1fda698;
      src10 <= 32'h4c6e6fbb;
      src11 <= 32'ha100ed14;
      src12 <= 32'h27fe1b4b;
      src13 <= 32'h78aff58e;
      src14 <= 32'had9d1f42;
      src15 <= 32'hc3121af6;
      src16 <= 32'hfbe86a8e;
      src17 <= 32'h1eeed219;
      src18 <= 32'ha614be3;
      src19 <= 32'h41aef3f7;
      src20 <= 32'h656fa7e6;
      src21 <= 32'h40aaec7a;
      src22 <= 32'he8a56f31;
      src23 <= 32'h986cc8d5;
      src24 <= 32'h9135087;
      src25 <= 32'hcad00273;
      src26 <= 32'h57030ede;
      src27 <= 32'h29deb984;
      src28 <= 32'h4a294067;
      src29 <= 32'h8513d91e;
      src30 <= 32'ha08c3a00;
      src31 <= 32'h88083ebc;
   end
endmodule

